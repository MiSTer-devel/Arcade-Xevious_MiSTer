library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity terrain_2a is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of terrain_2a is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"20",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"03",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"00",X"20",X"40",X"11",X"11",X"15",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"16",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"00",X"00",X"02",X"54",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"41",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"60",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",
		X"04",X"00",X"00",X"00",X"60",X"40",X"05",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"33",X"20",X"22",X"22",X"22",X"22",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"26",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"02",X"06",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"20",X"22",X"22",X"06",X"00",X"00",X"00",X"00",X"00",
		X"04",X"40",X"00",X"00",X"00",X"40",X"30",X"73",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"51",X"00",X"22",X"22",X"20",X"02",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"22",X"62",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"20",X"22",X"22",X"02",X"06",X"00",X"00",X"64",X"00",
		X"04",X"40",X"00",X"00",X"06",X"02",X"04",X"00",X"00",X"40",X"02",X"00",X"06",X"00",X"00",X"00",
		X"06",X"51",X"40",X"00",X"00",X"00",X"06",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"04",X"00",X"00",X"20",X"00",
		X"07",X"00",X"02",X"60",X"00",X"02",X"04",X"00",X"00",X"24",X"04",X"60",X"00",X"00",X"00",X"00",
		X"00",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"06",X"01",
		X"07",X"00",X"22",X"60",X"06",X"20",X"40",X"00",X"40",X"42",X"02",X"00",X"00",X"00",X"00",X"00",
		X"06",X"50",X"00",X"00",X"00",X"07",X"13",X"01",X"00",X"00",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"10",
		X"00",X"40",X"00",X"00",X"00",X"00",X"40",X"00",X"22",X"24",X"00",X"00",X"00",X"00",X"00",X"00",
		X"30",X"50",X"00",X"00",X"51",X"00",X"00",X"10",X"66",X"00",X"00",X"26",X"22",X"22",X"22",X"22",
		X"22",X"24",X"22",X"22",X"62",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"10",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"24",X"40",X"02",X"00",X"00",X"00",X"00",X"00",X"40",
		X"34",X"50",X"00",X"70",X"00",X"00",X"00",X"00",X"10",X"60",X"00",X"20",X"22",X"22",X"22",X"22",
		X"22",X"22",X"22",X"22",X"02",X"66",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",
		X"40",X"40",X"00",X"00",X"00",X"00",X"02",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"32",X"05",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"23",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"26",X"22",X"22",X"22",X"22",X"22",X"22",X"12",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",
		X"40",X"40",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"64",
		X"50",X"05",X"50",X"05",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"22",X"22",X"22",X"22",X"22",X"02",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"06",
		X"40",X"46",X"00",X"00",X"00",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"03",X"05",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"02",X"06",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"33",X"17",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"63",X"06",X"00",X"00",X"20",
		X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"70",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"20",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"13",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"01",X"00",X"20",X"54",
		X"11",X"20",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"36",
		X"30",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"02",X"00",X"00",X"00",X"10",X"02",X"44",X"07",
		X"00",X"13",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"74",X"00",X"00",X"00",X"07",X"15",X"31",
		X"03",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"02",X"66",X"66",X"00",X"00",X"13",X"51",X"00",
		X"00",X"00",X"00",X"21",X"02",X"60",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"04",
		X"40",X"00",X"24",X"22",X"22",X"22",X"22",X"02",X"00",X"40",X"00",X"50",X"51",X"00",X"14",X"05",
		X"01",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"02",X"06",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"10",X"11",X"02",X"04",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"22",X"00",X"00",X"04",X"00",X"04",
		X"40",X"00",X"26",X"22",X"22",X"22",X"22",X"22",X"24",X"40",X"15",X"51",X"40",X"01",X"10",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"02",X"06",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"01",X"04",X"00",X"00",X"00",X"00",X"50",X"00",X"00",
		X"00",X"00",X"30",X"00",X"00",X"00",X"04",X"00",X"00",X"60",X"00",X"02",X"00",X"04",X"00",X"04",
		X"40",X"60",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"05",X"00",X"00",X"00",X"40",X"07",
		X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"66",X"66",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"30",X"01",X"06",X"00",X"00",X"00",X"00",X"05",X"00",
		X"00",X"00",X"10",X"01",X"02",X"00",X"06",X"00",X"00",X"06",X"00",X"00",X"20",X"40",X"00",X"04",
		X"40",X"40",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"05",X"00",X"00",X"00",X"00",X"27",X"37",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"02",X"20",X"00",X"00",X"11",X"42",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"11",X"06",X"40",X"00",X"20",X"60",X"00",X"00",X"00",X"00",X"02",X"24",X"24",
		X"60",X"44",X"00",X"00",X"00",X"00",X"10",X"05",X"00",X"00",X"00",X"00",X"10",X"27",X"02",X"11",
		X"00",X"00",X"00",X"04",X"04",X"40",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"22",X"22",X"00",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"24",X"06",X"50",X"11",X"11",X"05",X"20",X"22",X"22",
		X"60",X"42",X"00",X"00",X"00",X"10",X"05",X"00",X"00",X"00",X"00",X"60",X"20",X"02",X"10",X"00",
		X"11",X"51",X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"01",X"40",X"04",X"14",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"60",X"22",X"22",X"42",X"02",X"10",X"00",X"00",X"30",X"00",X"00",X"00",
		X"40",X"60",X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"60",X"40",X"20",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"40",X"00",X"40",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"25",X"04",X"00",X"00",X"01",X"00",
		X"00",X"00",X"00",X"00",X"00",X"22",X"02",X"24",X"00",X"70",X"00",X"00",X"00",X"10",X"01",X"00",
		X"40",X"04",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"20",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"07",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"64",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"30",X"10",
		X"40",X"04",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"04",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"42",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"00",X"03",X"20",X"20",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"10",X"00",
		X"77",X"42",X"00",X"00",X"07",X"00",X"00",X"00",X"40",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"04",X"00",X"40",X"00",X"00",X"00",X"00",X"33",X"00",X"20",X"04",X"70",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"42",X"02",X"00",X"00",X"70",X"07",X"00",X"00",X"00",X"10",X"00",
		X"71",X"60",X"06",X"00",X"00",X"00",X"40",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"07",X"20",X"00",X"04",X"03",X"00",X"00",
		X"00",X"00",X"00",X"00",X"20",X"04",X"00",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"00",X"03",
		X"01",X"07",X"00",X"12",X"00",X"00",X"04",X"02",X"24",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"20",X"42",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"07",X"00",X"00",X"50",
		X"10",X"70",X"00",X"10",X"00",X"00",X"20",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"57",X"00",X"30",
		X"00",X"01",X"07",X"03",X"06",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"66",X"00",X"00",X"00",X"30",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"22",X"22",X"22",X"22",X"16",X"00",X"00",
		X"13",X"11",X"70",X"01",X"20",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"40",X"00",X"00",X"00",X"00",X"05",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"30",X"71",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",
		X"00",X"10",X"10",X"17",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"24",X"00",X"00",X"10",X"00",X"00",
		X"00",X"50",X"00",X"71",X"05",X"10",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"20",X"22",X"00",X"00",X"10",X"00",X"00",
		X"00",X"70",X"00",X"01",X"37",X"37",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"22",X"36",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",
		X"00",X"00",X"00",X"10",X"71",X"13",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"22",X"44",X"10",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"00",
		X"30",X"07",X"00",X"00",X"51",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"22",X"44",X"00",X"10",X"00",X"00",
		X"00",X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"77",X"00",
		X"07",X"00",X"40",X"00",X"00",X"00",X"51",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"42",X"40",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"33",
		X"00",X"00",X"00",X"04",X"04",X"00",X"00",X"15",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"02",X"04",X"00",X"00",X"00",X"00",X"01",X"00",X"00",
		X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"40",X"40",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"06",X"20",X"26",X"04",X"00",X"00",X"00",X"00",X"03",X"00",X"00",
		X"00",X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"44",X"00",X"00",X"10",X"11",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"66",X"00",X"62",X"00",X"42",X"00",X"00",X"00",X"00",X"07",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"05",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"00",X"00",X"04",X"00",X"20",X"04",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"10",X"11",X"55",X"15",X"11",
		X"51",X"11",X"15",X"11",X"11",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"51",X"11",
		X"15",X"11",X"15",X"00",X"42",X"10",X"35",X"51",X"00",X"04",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"04",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"15",X"00",X"00",X"10",X"11",X"51",X"01",X"00",X"00",X"50",X"51",X"00",X"50",X"05",
		X"05",X"00",X"00",X"06",X"15",X"05",X"00",X"00",X"01",X"42",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"31",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"15",X"05",X"00",X"60",X"72",X"73",
		X"22",X"62",X"40",X"02",X"01",X"00",X"00",X"00",X"10",X"02",X"04",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"00",X"00",X"44",X"00",X"00",X"00",X"00",
		X"70",X"33",X"00",X"77",X"33",X"00",X"22",X"60",X"22",X"26",X"04",X"00",X"24",X"00",X"00",X"60",
		X"00",X"00",X"40",X"00",X"01",X"00",X"00",X"00",X"10",X"40",X"42",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"01",X"00",X"00",X"00",X"44",X"00",X"00",X"00",
		X"50",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"04",X"01",X"00",X"00",X"00",X"00",X"25",X"20",X"04",X"10",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"06",X"00",X"00",X"00",X"00",X"02",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"00",X"00",X"00",X"00",X"44",X"00",X"00",
		X"70",X"00",X"00",X"00",X"70",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"40",X"01",X"00",X"00",X"00",X"00",X"05",X"04",X"42",X"10",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"60",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"44",X"00",
		X"50",X"01",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"54",X"00",X"00",X"00",X"00",X"21",X"04",X"20",X"14",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"44",
		X"00",X"50",X"00",X"00",X"11",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"03",X"04",X"00",X"42",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"11",X"01",X"00",X"00",
		X"04",X"00",X"51",X"51",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"15",X"11",X"11",X"00",X"00",
		X"40",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"50",X"04",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"11",X"02",X"00",X"00",
		X"00",X"44",X"00",X"00",X"00",X"20",X"00",X"26",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"14",X"00",X"00",X"00",X"00",X"50",X"02",X"00",X"75",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"22",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"02",X"02",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"16",X"00",X"00",X"00",X"00",X"50",X"40",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"22",X"22",
		X"02",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"20",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"70",X"00",X"00",X"00",X"00",X"50",X"02",X"66",X"07",X"00",X"00",X"00",
		X"00",X"00",X"05",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"20",X"02",X"20",
		X"22",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"00",X"22",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"60",X"01",X"00",X"00",X"00",X"00",X"30",X"20",X"06",X"00",X"00",X"00",X"00",
		X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"02",X"00",X"22",X"00",X"00",
		X"22",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"02",X"00",X"00",X"00",
		X"00",X"00",X"40",X"54",X"05",X"00",X"00",X"00",X"00",X"00",X"45",X"01",X"00",X"00",X"00",X"00",
		X"00",X"00",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"00",X"00",X"00",X"22",X"02",X"00",
		X"00",X"40",X"06",X"55",X"00",X"00",X"00",X"00",X"00",X"00",X"05",X"54",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
