library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity xevious_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(13 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of xevious_cpu1 is
	type rom is array(0 to  16383) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"3E",X"10",X"32",X"00",X"71",X"C3",X"2E",X"01",X"87",X"D2",X"4F",X"00",X"25",X"C3",X"4F",X"00",
		X"A7",X"F2",X"4F",X"00",X"25",X"C3",X"4F",X"00",X"A7",X"F0",X"ED",X"44",X"C9",X"33",X"33",X"C9",
		X"06",X"03",X"21",X"80",X"81",X"AF",X"18",X"2C",X"EB",X"CD",X"28",X"01",X"29",X"29",X"19",X"C9",
		X"E1",X"DD",X"75",X"00",X"DD",X"74",X"01",X"C9",X"E5",X"D5",X"C5",X"F5",X"32",X"30",X"68",X"21",
		X"20",X"68",X"36",X"00",X"36",X"01",X"CD",X"96",X"00",X"F1",X"C1",X"D1",X"E1",X"FB",X"C9",X"85",
		X"6F",X"D0",X"24",X"C9",X"1A",X"8E",X"27",X"77",X"13",X"23",X"10",X"F8",X"DC",X"09",X"13",X"CD",
		X"11",X"13",X"C3",X"3A",X"13",X"FF",X"D9",X"ED",X"A0",X"EA",X"93",X"00",X"08",X"3E",X"10",X"32",
		X"00",X"71",X"2A",X"04",X"80",X"7E",X"A7",X"28",X"19",X"36",X"00",X"2C",X"2C",X"4E",X"2C",X"46",
		X"2C",X"5E",X"2C",X"56",X"2C",X"D5",X"5E",X"2C",X"56",X"2C",X"22",X"04",X"80",X"EB",X"D1",X"32",
		X"00",X"71",X"08",X"D9",X"ED",X"45",X"21",X"00",X"82",X"11",X"80",X"87",X"01",X"40",X"00",X"ED",
		X"B0",X"21",X"00",X"83",X"11",X"80",X"97",X"01",X"40",X"00",X"ED",X"B0",X"21",X"00",X"81",X"11",
		X"80",X"A7",X"01",X"40",X"00",X"ED",X"B0",X"2A",X"20",X"80",X"7D",X"A4",X"32",X"03",X"80",X"32",
		X"70",X"D0",X"3A",X"AD",X"85",X"A7",X"28",X"12",X"3A",X"18",X"80",X"FE",X"BB",X"28",X"FE",X"CD",
		X"15",X"01",X"CB",X"7D",X"C8",X"3E",X"01",X"32",X"02",X"80",X"3E",X"01",X"32",X"00",X"80",X"21",
		X"18",X"80",X"01",X"03",X"71",X"11",X"00",X"70",X"EB",X"3A",X"00",X"71",X"E6",X"E0",X"78",X"06",
		X"00",X"20",X"05",X"D9",X"32",X"00",X"71",X"C9",X"E5",X"2A",X"06",X"80",X"77",X"2C",X"2C",X"71",
		X"2C",X"70",X"2C",X"73",X"2C",X"72",X"2C",X"D1",X"73",X"2C",X"72",X"2C",X"22",X"06",X"80",X"C9",
		X"11",X"00",X"70",X"18",X"D4",X"11",X"00",X"68",X"06",X"08",X"1A",X"1F",X"CB",X"1D",X"1F",X"CB",
		X"1C",X"13",X"10",X"F6",X"22",X"16",X"80",X"C9",X"21",X"00",X"00",X"C3",X"08",X"00",X"F3",X"ED",
		X"56",X"AF",X"32",X"30",X"68",X"32",X"0A",X"80",X"32",X"10",X"D0",X"32",X"30",X"D0",X"32",X"20",
		X"68",X"32",X"21",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"01",X"20",X"00",X"21",X"00",X"68",
		X"70",X"23",X"0D",X"20",X"FB",X"31",X"00",X"D0",X"06",X"00",X"58",X"FD",X"21",X"3D",X"03",X"DD",
		X"21",X"31",X"03",X"21",X"00",X"00",X"DD",X"56",X"00",X"DD",X"4E",X"01",X"15",X"28",X"2D",X"FD",
		X"35",X"00",X"20",X"0E",X"32",X"30",X"68",X"78",X"86",X"12",X"23",X"13",X"79",X"BA",X"20",X"F4",
		X"18",X"14",X"EB",X"32",X"30",X"68",X"1A",X"80",X"BE",X"20",X"1E",X"23",X"13",X"79",X"BC",X"20",
		X"F2",X"EB",X"FE",X"CF",X"28",X"0A",X"DD",X"23",X"DD",X"23",X"18",X"CA",X"FD",X"23",X"18",X"BF",
		X"78",X"C6",X"11",X"38",X"0D",X"47",X"C3",X"5B",X"01",X"7C",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",
		X"CB",X"3F",X"32",X"00",X"85",X"AF",X"32",X"AD",X"85",X"CD",X"67",X"03",X"11",X"3E",X"03",X"32",
		X"30",X"68",X"13",X"1A",X"6F",X"13",X"1A",X"67",X"A7",X"28",X"0D",X"13",X"1A",X"A7",X"28",X"EF",
		X"77",X"13",X"01",X"C0",X"FF",X"09",X"18",X"F4",X"3A",X"00",X"85",X"FE",X"10",X"28",X"08",X"32",
		X"CF",X"C4",X"32",X"30",X"68",X"18",X"FB",X"3E",X"18",X"32",X"CF",X"C4",X"3E",X"14",X"32",X"8F",
		X"C4",X"31",X"80",X"A7",X"AF",X"21",X"00",X"80",X"11",X"01",X"80",X"01",X"FF",X"03",X"77",X"ED",
		X"B0",X"32",X"30",X"68",X"21",X"80",X"87",X"77",X"2C",X"20",X"FC",X"21",X"80",X"97",X"77",X"2C",
		X"20",X"FC",X"21",X"80",X"A7",X"77",X"2C",X"20",X"FC",X"32",X"AD",X"85",X"21",X"00",X"92",X"22",
		X"04",X"80",X"22",X"06",X"80",X"77",X"2C",X"20",X"FC",X"3E",X"01",X"32",X"20",X"68",X"32",X"22",
		X"68",X"32",X"23",X"68",X"21",X"55",X"03",X"01",X"06",X"A1",X"CD",X"10",X"01",X"FB",X"11",X"74",
		X"85",X"21",X"00",X"00",X"0E",X"10",X"06",X"00",X"78",X"86",X"12",X"23",X"47",X"79",X"BC",X"20",
		X"F7",X"13",X"79",X"C6",X"10",X"4F",X"FE",X"50",X"20",X"EC",X"06",X"07",X"21",X"71",X"85",X"7E",
		X"A7",X"20",X"15",X"23",X"05",X"20",X"F8",X"3E",X"18",X"32",X"D1",X"C4",X"3E",X"14",X"32",X"91",
		X"C4",X"3E",X"0F",X"32",X"AC",X"85",X"18",X"06",X"78",X"32",X"D1",X"C4",X"18",X"FE",X"16",X"08",
		X"21",X"00",X"68",X"DD",X"21",X"D5",X"C4",X"FD",X"21",X"95",X"C4",X"01",X"00",X"00",X"7E",X"1F",
		X"3F",X"CB",X"11",X"1F",X"3F",X"CB",X"10",X"DD",X"70",X"00",X"FD",X"71",X"00",X"DD",X"23",X"FD",
		X"23",X"23",X"15",X"20",X"E6",X"3A",X"AC",X"85",X"32",X"D3",X"C4",X"3A",X"18",X"80",X"87",X"38",
		X"26",X"FE",X"FE",X"20",X"07",X"3A",X"19",X"80",X"3C",X"CA",X"7E",X"02",X"3A",X"AC",X"85",X"3C",
		X"FE",X"10",X"20",X"01",X"AF",X"32",X"AC",X"85",X"32",X"D3",X"C4",X"26",X"A0",X"6F",X"3E",X"01",
		X"77",X"CD",X"5B",X"03",X"C3",X"7E",X"02",X"CD",X"67",X"03",X"3E",X"27",X"0E",X"18",X"21",X"C4",
		X"C6",X"06",X"22",X"E5",X"D1",X"12",X"13",X"05",X"20",X"FB",X"06",X"40",X"2B",X"05",X"20",X"FC",
		X"0D",X"20",X"EE",X"21",X"C5",X"B6",X"3E",X"64",X"CD",X"1B",X"03",X"21",X"84",X"B6",X"3E",X"A4",
		X"CD",X"1B",X"03",X"21",X"85",X"B6",X"3E",X"E4",X"CD",X"1B",X"03",X"CD",X"5B",X"03",X"3A",X"18",
		X"80",X"CB",X"7F",X"28",X"F9",X"CD",X"5B",X"03",X"C3",X"88",X"03",X"0E",X"0C",X"E5",X"D1",X"06",
		X"11",X"12",X"13",X"13",X"05",X"20",X"FA",X"06",X"80",X"2B",X"05",X"20",X"FC",X"0D",X"20",X"ED",
		X"C9",X"79",X"80",X"83",X"88",X"91",X"92",X"95",X"97",X"A1",X"A8",X"B1",X"CF",X"01",X"00",X"CF",
		X"C5",X"1B",X"0A",X"16",X"00",X"D1",X"C5",X"1B",X"18",X"16",X"00",X"53",X"C6",X"1C",X"18",X"1E",
		X"17",X"0D",X"00",X"00",X"00",X"05",X"05",X"05",X"05",X"05",X"05",X"E5",X"21",X"00",X"00",X"2D",
		X"20",X"FD",X"25",X"20",X"FA",X"E1",X"C9",X"21",X"80",X"97",X"01",X"98",X"24",X"CD",X"7D",X"03",
		X"21",X"00",X"78",X"0E",X"80",X"CD",X"7D",X"03",X"21",X"00",X"B0",X"0E",X"CF",X"32",X"30",X"68",
		X"78",X"77",X"23",X"7C",X"B9",X"20",X"F6",X"C9",X"21",X"D2",X"03",X"11",X"60",X"85",X"01",X"08",
		X"00",X"ED",X"B0",X"16",X"08",X"21",X"00",X"68",X"7E",X"1F",X"CB",X"19",X"1F",X"CB",X"18",X"23",
		X"15",X"20",X"F5",X"21",X"CA",X"03",X"78",X"E6",X"03",X"CB",X"27",X"85",X"6F",X"7E",X"32",X"63",
		X"85",X"23",X"7E",X"32",X"64",X"85",X"21",X"CA",X"03",X"79",X"1F",X"E6",X"06",X"85",X"6F",X"7E",
		X"32",X"65",X"85",X"23",X"7E",X"32",X"66",X"85",X"18",X"10",X"02",X"03",X"02",X"01",X"01",X"02",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"02",X"02",X"F3",X"3E",X"10",X"32",X"00",X"71",
		X"AF",X"32",X"30",X"68",X"32",X"0A",X"80",X"32",X"10",X"D0",X"32",X"30",X"D0",X"32",X"20",X"68",
		X"32",X"21",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"21",X"00",X"80",X"11",X"01",X"80",X"01",
		X"FF",X"01",X"36",X"00",X"ED",X"B0",X"21",X"00",X"92",X"22",X"04",X"80",X"22",X"06",X"80",X"36",
		X"00",X"2C",X"20",X"FB",X"21",X"5B",X"04",X"11",X"80",X"82",X"01",X"40",X"00",X"ED",X"B0",X"3E",
		X"01",X"32",X"20",X"68",X"32",X"22",X"68",X"32",X"23",X"68",X"32",X"AD",X"85",X"21",X"60",X"85",
		X"01",X"08",X"A1",X"CD",X"10",X"01",X"FB",X"2A",X"00",X"80",X"2D",X"20",X"FA",X"24",X"22",X"00",
		X"80",X"DD",X"21",X"80",X"82",X"06",X"20",X"C5",X"CD",X"54",X"04",X"C1",X"DD",X"23",X"DD",X"23",
		X"10",X"F5",X"18",X"E3",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"E9",X"9B",X"04",X"BB",X"14",X"00",
		X"30",X"D0",X"33",X"B3",X"33",X"E5",X"33",X"08",X"0F",X"9E",X"3B",X"E3",X"3B",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",
		X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"27",X"17",X"62",X"18",X"CD",X"E1",X"06",X"CD",X"0D",
		X"07",X"CD",X"2A",X"07",X"CD",X"D9",X"10",X"3A",X"17",X"80",X"07",X"2F",X"E6",X"01",X"32",X"20",
		X"80",X"3E",X"01",X"32",X"2A",X"80",X"3E",X"F8",X"32",X"14",X"80",X"21",X"0E",X"0C",X"01",X"02",
		X"61",X"F3",X"CD",X"10",X"01",X"FB",X"AF",X"32",X"23",X"80",X"3A",X"29",X"80",X"A7",X"20",X"1B",
		X"3E",X"02",X"32",X"28",X"80",X"F7",X"3A",X"28",X"80",X"3D",X"21",X"40",X"0C",X"CF",X"5E",X"23",
		X"56",X"EB",X"E9",X"CD",X"81",X"08",X"3A",X"29",X"80",X"A7",X"C8",X"CD",X"F0",X"06",X"AF",X"32",
		X"28",X"80",X"3C",X"32",X"2A",X"80",X"CD",X"0D",X"07",X"CD",X"2A",X"07",X"CD",X"3C",X"08",X"CD",
		X"D5",X"0D",X"CD",X"DC",X"07",X"CD",X"AA",X"08",X"F7",X"CD",X"01",X"08",X"CD",X"23",X"08",X"3A",
		X"1B",X"80",X"A7",X"C8",X"32",X"23",X"80",X"AF",X"32",X"21",X"80",X"32",X"1B",X"80",X"21",X"80",
		X"81",X"77",X"2C",X"77",X"2C",X"77",X"2C",X"EB",X"21",X"0A",X"0C",X"3A",X"17",X"80",X"07",X"07",
		X"07",X"E6",X"03",X"D7",X"7E",X"EB",X"77",X"2C",X"2C",X"2C",X"2C",X"36",X"00",X"2C",X"36",X"00",
		X"2C",X"EB",X"3A",X"17",X"80",X"07",X"07",X"07",X"E6",X"03",X"EE",X"03",X"28",X"02",X"3E",X"01",
		X"21",X"10",X"0C",X"CF",X"4E",X"23",X"7E",X"67",X"69",X"3A",X"17",X"80",X"2F",X"0F",X"0F",X"E6",
		X"07",X"CF",X"EB",X"1A",X"77",X"2C",X"13",X"1A",X"77",X"2C",X"36",X"01",X"2C",X"3A",X"17",X"80",
		X"2F",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"3E",X"00",X"20",X"01",X"3C",X"77",X"3A",X"22",X"80",
		X"A7",X"28",X"10",X"21",X"80",X"81",X"11",X"C0",X"81",X"01",X"40",X"00",X"ED",X"B0",X"3E",X"01",
		X"32",X"01",X"A0",X"21",X"83",X"81",X"35",X"3A",X"87",X"81",X"4F",X"21",X"B3",X"3E",X"D7",X"7E",
		X"32",X"13",X"80",X"21",X"00",X"0D",X"22",X"10",X"80",X"79",X"21",X"00",X"A4",X"CF",X"7E",X"32",
		X"85",X"81",X"23",X"7E",X"32",X"86",X"81",X"AF",X"32",X"2B",X"80",X"32",X"2C",X"80",X"32",X"2D",
		X"80",X"32",X"22",X"84",X"32",X"44",X"80",X"CD",X"0D",X"07",X"CD",X"47",X"07",X"CD",X"D5",X"0D",
		X"CD",X"68",X"0F",X"21",X"62",X"18",X"22",X"BE",X"82",X"21",X"BB",X"14",X"22",X"82",X"82",X"AF",
		X"32",X"2A",X"80",X"3C",X"32",X"01",X"A0",X"3E",X"A0",X"32",X"41",X"80",X"CD",X"7F",X"07",X"F7",
		X"21",X"41",X"80",X"35",X"C0",X"CD",X"B7",X"07",X"F7",X"3A",X"2A",X"80",X"A7",X"C8",X"CD",X"47",
		X"07",X"3E",X"40",X"32",X"41",X"80",X"3A",X"11",X"80",X"D6",X"0E",X"FE",X"36",X"30",X"0B",X"21",
		X"87",X"81",X"34",X"3E",X"10",X"BE",X"20",X"02",X"36",X"06",X"3A",X"16",X"80",X"2F",X"07",X"07",
		X"07",X"E6",X"03",X"21",X"34",X"0C",X"D7",X"4E",X"3A",X"88",X"81",X"91",X"30",X"01",X"AF",X"32",
		X"88",X"81",X"F7",X"21",X"41",X"80",X"35",X"C0",X"21",X"40",X"79",X"11",X"41",X"79",X"01",X"0D",
		X"00",X"36",X"00",X"ED",X"B0",X"3A",X"83",X"81",X"A7",X"20",X"37",X"C3",X"43",X"11",X"3A",X"22",
		X"80",X"A7",X"28",X"1A",X"CD",X"0D",X"07",X"CD",X"47",X"07",X"CD",X"D5",X"0D",X"CD",X"6A",X"08",
		X"3E",X"80",X"32",X"41",X"80",X"F7",X"21",X"41",X"80",X"35",X"C0",X"CD",X"49",X"08",X"3A",X"C3",
		X"81",X"A7",X"28",X"17",X"CD",X"6D",X"07",X"3A",X"21",X"80",X"EE",X"01",X"32",X"21",X"80",X"C3",
		X"93",X"05",X"3A",X"C3",X"81",X"A7",X"20",X"EC",X"C3",X"93",X"05",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"D5",X"0D",X"CD",X"5D",X"08",X"3E",X"80",X"32",X"41",X"80",X"F7",X"21",X"41",X"80",
		X"35",X"C0",X"CD",X"49",X"08",X"3A",X"21",X"80",X"A7",X"CA",X"BB",X"04",X"CD",X"6D",X"07",X"AF",
		X"32",X"21",X"80",X"C3",X"BB",X"04",X"21",X"00",X"78",X"11",X"00",X"10",X"36",X"00",X"23",X"1B",
		X"7B",X"B2",X"20",X"F8",X"21",X"00",X"90",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",
		X"20",X"F8",X"21",X"00",X"A0",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",
		X"C9",X"21",X"00",X"78",X"11",X"00",X"08",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",
		X"21",X"00",X"79",X"11",X"40",X"00",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"74",
		X"79",X"11",X"06",X"00",X"36",X"00",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B0",
		X"11",X"00",X"08",X"36",X"24",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C0",X"11",X"00",
		X"08",X"36",X"24",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B8",X"11",X"00",X"08",
		X"36",X"03",X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C8",X"11",X"00",X"08",X"36",X"00",
		X"23",X"1B",X"7B",X"B2",X"20",X"F8",X"C9",X"21",X"00",X"B8",X"11",X"00",X"08",X"36",X"00",X"23",
		X"1B",X"7B",X"B2",X"20",X"F8",X"21",X"00",X"C8",X"3E",X"88",X"06",X"1C",X"77",X"23",X"3C",X"10",
		X"FB",X"21",X"00",X"C8",X"11",X"1C",X"C8",X"01",X"E4",X"07",X"ED",X"B0",X"C9",X"06",X"40",X"21",
		X"80",X"81",X"11",X"C0",X"81",X"4E",X"1A",X"77",X"79",X"12",X"2C",X"1C",X"10",X"F7",X"C9",X"3A",
		X"21",X"80",X"21",X"E5",X"0B",X"CF",X"5E",X"23",X"56",X"21",X"17",X"12",X"06",X"0A",X"0E",X"C0",
		X"CD",X"1F",X"14",X"21",X"19",X"10",X"11",X"DF",X"0B",X"06",X"06",X"0E",X"C0",X"CD",X"1F",X"14",
		X"11",X"FD",X"0B",X"21",X"1B",X"13",X"06",X"0D",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"1B",X"15",
		X"3A",X"83",X"81",X"CD",X"4F",X"14",X"C9",X"21",X"17",X"12",X"06",X"0A",X"3E",X"24",X"0E",X"C0",
		X"CD",X"5D",X"14",X"21",X"19",X"10",X"06",X"06",X"3E",X"24",X"0E",X"C0",X"CD",X"5D",X"14",X"06",
		X"10",X"21",X"1B",X"15",X"3E",X"24",X"0E",X"C0",X"CD",X"5D",X"14",X"C9",X"21",X"1F",X"16",X"11",
		X"CD",X"3E",X"06",X"13",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"21",X"10",X"11",X"E0",X"3E",X"06",
		X"07",X"CD",X"1F",X"14",X"21",X"21",X"10",X"06",X"07",X"0E",X"B0",X"3E",X"1A",X"CD",X"5D",X"14",
		X"C9",X"21",X"23",X"09",X"11",X"D9",X"0B",X"06",X"06",X"0E",X"C0",X"CD",X"1F",X"14",X"25",X"3A",
		X"29",X"80",X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"CD",X"4F",X"14",X"3A",X"29",X"80",X"E6",X"0F",
		X"C3",X"4F",X"14",X"3A",X"29",X"80",X"FE",X"01",X"28",X"01",X"AF",X"21",X"B1",X"0B",X"CF",X"5E",
		X"23",X"56",X"21",X"19",X"15",X"06",X"12",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"17",X"15",X"11",
		X"A0",X"0B",X"06",X"11",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"18",X"11",X"06",X"09",X"0E",X"C0",
		X"3E",X"24",X"CD",X"5D",X"14",X"21",X"1A",X"12",X"06",X"0A",X"C3",X"5D",X"14",X"21",X"18",X"11",
		X"11",X"97",X"0B",X"06",X"09",X"0E",X"C0",X"C3",X"1F",X"14",X"CD",X"5D",X"08",X"3A",X"21",X"80",
		X"21",X"E5",X"0B",X"CF",X"5E",X"23",X"56",X"21",X"1A",X"12",X"06",X"0A",X"0E",X"C0",X"C3",X"1F",
		X"14",X"3A",X"01",X"80",X"4F",X"E6",X"0F",X"C0",X"79",X"0F",X"0F",X"0F",X"0F",X"E6",X"01",X"28",
		X"0D",X"21",X"1C",X"12",X"11",X"8C",X"0B",X"06",X"0B",X"0E",X"C0",X"C3",X"1F",X"14",X"21",X"1C",
		X"12",X"06",X"0B",X"0E",X"C0",X"3E",X"24",X"C3",X"5D",X"14",X"21",X"04",X"00",X"22",X"0C",X"80",
		X"0E",X"C8",X"21",X"09",X"15",X"11",X"9F",X"0A",X"06",X"12",X"CD",X"1F",X"14",X"21",X"0A",X"16",
		X"11",X"B1",X"0A",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0B",X"15",X"11",X"C4",X"0A",X"06",X"12",
		X"CD",X"1F",X"14",X"21",X"0C",X"16",X"11",X"D6",X"0A",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0D",
		X"17",X"11",X"E9",X"0A",X"06",X"14",X"CD",X"1F",X"14",X"21",X"0E",X"17",X"11",X"FD",X"0A",X"06",
		X"13",X"CD",X"1F",X"14",X"21",X"0F",X"17",X"11",X"10",X"0B",X"06",X"11",X"CD",X"1F",X"14",X"21",
		X"10",X"15",X"3E",X"F9",X"CD",X"4F",X"14",X"0E",X"B8",X"21",X"09",X"15",X"3E",X"0D",X"06",X"12",
		X"CD",X"5D",X"14",X"21",X"0A",X"16",X"3E",X"0D",X"06",X"13",X"CD",X"5D",X"14",X"21",X"0B",X"15",
		X"3E",X"11",X"06",X"02",X"CD",X"5D",X"14",X"3E",X"15",X"06",X"0F",X"CD",X"5D",X"14",X"3E",X"11",
		X"CD",X"4F",X"14",X"21",X"0C",X"16",X"3E",X"13",X"06",X"02",X"CD",X"5D",X"14",X"3E",X"17",X"06",
		X"10",X"CD",X"5D",X"14",X"3E",X"13",X"CD",X"4F",X"14",X"21",X"0D",X"17",X"3E",X"13",X"06",X"02",
		X"CD",X"5D",X"14",X"3E",X"17",X"06",X"10",X"CD",X"5D",X"14",X"3E",X"0F",X"CD",X"4F",X"14",X"3E",
		X"13",X"CD",X"4F",X"14",X"21",X"0E",X"17",X"3E",X"13",X"CD",X"4F",X"14",X"3E",X"19",X"06",X"11",
		X"CD",X"5D",X"14",X"3E",X"18",X"CD",X"4F",X"14",X"21",X"0F",X"17",X"3E",X"18",X"06",X"02",X"CD",
		X"5D",X"14",X"3E",X"19",X"CD",X"4F",X"14",X"3E",X"18",X"06",X"0E",X"CD",X"5D",X"14",X"21",X"10",
		X"15",X"3E",X"18",X"CD",X"4F",X"14",X"0E",X"C0",X"21",X"0B",X"15",X"11",X"60",X"0A",X"06",X"11",
		X"CD",X"1F",X"14",X"21",X"0C",X"13",X"11",X"71",X"0A",X"06",X"0E",X"CD",X"1F",X"14",X"21",X"0D",
		X"14",X"11",X"7F",X"0A",X"06",X"10",X"CD",X"1F",X"14",X"21",X"0E",X"15",X"11",X"8F",X"0A",X"06",
		X"10",X"CD",X"1F",X"14",X"3E",X"1A",X"0E",X"B0",X"21",X"0B",X"15",X"06",X"11",X"CD",X"5D",X"14",
		X"21",X"0C",X"13",X"06",X"0E",X"CD",X"5D",X"14",X"21",X"0D",X"14",X"06",X"10",X"CD",X"5D",X"14",
		X"21",X"0E",X"15",X"06",X"10",X"C3",X"5D",X"14",X"21",X"0A",X"16",X"11",X"21",X"0B",X"0E",X"C0",
		X"06",X"13",X"CD",X"1F",X"14",X"21",X"0B",X"15",X"11",X"34",X"0B",X"06",X"12",X"CD",X"1F",X"14",
		X"21",X"0C",X"15",X"11",X"46",X"0B",X"06",X"12",X"CD",X"1F",X"14",X"21",X"0D",X"16",X"11",X"58",
		X"0B",X"06",X"13",X"CD",X"1F",X"14",X"21",X"0E",X"17",X"11",X"6B",X"0B",X"06",X"14",X"CD",X"1F",
		X"14",X"21",X"0F",X"17",X"11",X"7F",X"0B",X"06",X"0D",X"CD",X"1F",X"14",X"3E",X"1B",X"21",X"0A",
		X"16",X"0E",X"B0",X"06",X"13",X"CD",X"5D",X"14",X"21",X"0B",X"15",X"06",X"12",X"CD",X"5D",X"14",
		X"21",X"0C",X"15",X"06",X"12",X"CD",X"5D",X"14",X"21",X"0D",X"16",X"06",X"13",X"CD",X"5D",X"14",
		X"21",X"0E",X"17",X"06",X"14",X"CD",X"5D",X"14",X"21",X"0F",X"17",X"06",X"0D",X"C3",X"5D",X"14",
		X"2A",X"51",X"52",X"53",X"52",X"54",X"55",X"56",X"24",X"57",X"58",X"59",X"5A",X"5B",X"5C",X"5D",
		X"52",X"5E",X"5F",X"2A",X"60",X"61",X"62",X"63",X"64",X"65",X"66",X"67",X"68",X"69",X"6A",X"6B",
		X"6C",X"6D",X"6E",X"6F",X"70",X"71",X"72",X"73",X"74",X"75",X"76",X"77",X"78",X"79",X"7A",X"7B",
		X"7C",X"7D",X"7E",X"7F",X"80",X"81",X"82",X"83",X"84",X"85",X"86",X"87",X"7F",X"88",X"89",X"C0",
		X"C1",X"C2",X"C3",X"C2",X"C4",X"C5",X"C1",X"C6",X"C7",X"C1",X"C8",X"C1",X"C9",X"CA",X"CB",X"CA",
		X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"D3",X"D4",X"D5",X"D6",X"D7",X"D8",X"D9",X"DA",X"DB",
		X"DC",X"DD",X"DE",X"DF",X"E0",X"E1",X"E2",X"E3",X"E4",X"E5",X"E6",X"E7",X"E8",X"E9",X"EA",X"EB",
		X"EC",X"ED",X"EE",X"EF",X"F0",X"F1",X"F2",X"F3",X"F4",X"F5",X"F6",X"F7",X"F8",X"F9",X"FA",X"FB",
		X"FC",X"FD",X"FE",X"FF",X"A0",X"A1",X"A2",X"A3",X"A4",X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",
		X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",X"B5",X"B6",X"B7",X"B8",X"B9",X"BA",X"BB",
		X"BB",X"BB",X"BB",X"BB",X"BB",X"BC",X"BD",X"BD",X"BD",X"BE",X"BB",X"BB",X"BB",X"BB",X"BF",X"F0",
		X"F1",X"F2",X"BB",X"F3",X"F4",X"F4",X"F4",X"F4",X"F5",X"F6",X"F6",X"F6",X"F7",X"F4",X"F4",X"F4",
		X"F8",X"8A",X"8B",X"8C",X"8D",X"8E",X"8D",X"8F",X"90",X"87",X"91",X"92",X"93",X"94",X"87",X"95",
		X"96",X"97",X"98",X"99",X"9A",X"9B",X"9C",X"9D",X"9C",X"9E",X"9F",X"A0",X"A1",X"A2",X"A3",X"A4",
		X"A5",X"A6",X"A7",X"A8",X"A9",X"AA",X"AB",X"AC",X"AD",X"AE",X"AF",X"B0",X"B1",X"B2",X"B3",X"B4",
		X"B5",X"B6",X"B7",X"B8",X"A7",X"B9",X"9A",X"BA",X"AB",X"BB",X"AA",X"9A",X"BC",X"BD",X"BE",X"BF",
		X"C0",X"C1",X"C2",X"9A",X"C3",X"AA",X"C4",X"C5",X"C6",X"C7",X"C8",X"AB",X"BB",X"C9",X"CA",X"CA",
		X"CB",X"CC",X"CD",X"CE",X"CF",X"D0",X"D1",X"D2",X"CB",X"CA",X"CA",X"D3",X"D4",X"D5",X"D6",X"D7",
		X"AA",X"24",X"24",X"24",X"24",X"24",X"24",X"D8",X"D9",X"D9",X"D9",X"DA",X"12",X"17",X"1C",X"0E",
		X"1B",X"1D",X"24",X"0C",X"18",X"12",X"17",X"10",X"0A",X"16",X"0E",X"24",X"18",X"1F",X"0E",X"1B",
		X"19",X"1E",X"1C",X"11",X"24",X"1C",X"1D",X"0A",X"1B",X"1D",X"24",X"0B",X"1E",X"1D",X"1D",X"18",
		X"17",X"C7",X"0B",X"B5",X"0B",X"24",X"18",X"17",X"0E",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",
		X"24",X"18",X"17",X"15",X"22",X"24",X"24",X"18",X"17",X"0E",X"24",X"18",X"1B",X"24",X"1D",X"20",
		X"18",X"24",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"1C",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"1B",
		X"0E",X"0A",X"0D",X"22",X"2C",X"E9",X"0B",X"F3",X"0B",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",
		X"18",X"17",X"0E",X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"1D",X"20",X"18",X"1C",X"18",X"15",
		X"1F",X"0A",X"15",X"18",X"1E",X"24",X"15",X"0E",X"0F",X"1D",X"05",X"02",X"01",X"03",X"02",X"02",
		X"14",X"0C",X"24",X"0C",X"20",X"00",X"10",X"00",X"20",X"00",X"20",X"00",X"20",X"00",X"30",X"00",
		X"20",X"00",X"FF",X"FF",X"20",X"00",X"10",X"00",X"10",X"00",X"20",X"00",X"20",X"00",X"20",X"00",
		X"20",X"00",X"FF",X"FF",X"10",X"18",X"08",X"00",X"1A",X"17",X"18",X"07",X"3A",X"1B",X"1F",X"15",
		X"35",X"0D",X"48",X"0C",X"35",X"0D",X"A2",X"0D",X"CD",X"2A",X"07",X"CD",X"0D",X"07",X"CD",X"DC",
		X"07",X"CD",X"D5",X"0D",X"CD",X"AA",X"08",X"3E",X"40",X"32",X"41",X"80",X"11",X"65",X"0C",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"21",X"41",X"80",X"35",X"28",X"03",X"C3",X"E3",X"04",X"21",X"60",
		X"0D",X"22",X"1E",X"7A",X"21",X"60",X"16",X"22",X"1E",X"7B",X"21",X"30",X"0F",X"22",X"1E",X"7C",
		X"21",X"02",X"80",X"22",X"1E",X"79",X"AF",X"32",X"1E",X"7D",X"11",X"93",X"0C",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"1E",X"7D",X"3C",X"32",X"1E",X"7D",X"FE",X"10",X"28",X"0B",X"0F",X"E6",
		X"07",X"C6",X"30",X"32",X"1E",X"7C",X"C3",X"E3",X"04",X"3E",X"78",X"32",X"1E",X"7D",X"11",X"B7",
		X"0C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"1E",X"7D",X"3C",X"32",X"1E",X"7D",X"28",X"13",
		X"E6",X"07",X"C6",X"38",X"32",X"1E",X"7C",X"2A",X"1E",X"7B",X"3E",X"F0",X"CF",X"22",X"1E",X"7B",
		X"C3",X"E3",X"04",X"3E",X"10",X"32",X"1E",X"7D",X"11",X"E1",X"0C",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"3A",X"1E",X"7D",X"3D",X"32",X"1E",X"7D",X"28",X"0B",X"0F",X"E6",X"07",X"C6",X"30",X"32",
		X"1E",X"7C",X"C3",X"E3",X"04",X"AF",X"32",X"41",X"80",X"32",X"1E",X"79",X"11",X"05",X"0D",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",X"80",X"E6",X"01",X"C2",X"E3",X"04",X"21",X"41",X"80",
		X"35",X"28",X"0E",X"7E",X"E6",X"07",X"21",X"38",X"0C",X"D7",X"7E",X"CD",X"C6",X"09",X"C3",X"E3",
		X"04",X"CD",X"F0",X"06",X"3E",X"03",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"C3",X"E3",X"04",X"AF",X"32",X"21",X"80",X"32",X"87",X"81",X"32",X"88",X"81",X"21",
		X"B3",X"3E",X"D7",X"7E",X"32",X"13",X"80",X"21",X"00",X"0D",X"22",X"10",X"80",X"AF",X"21",X"00",
		X"A4",X"CF",X"7E",X"32",X"85",X"81",X"23",X"7E",X"32",X"86",X"81",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"D5",X"0D",X"CD",X"DC",X"07",X"CD",X"E8",X"09",X"AF",X"32",X"2B",X"80",X"32",X"2C",
		X"80",X"32",X"2D",X"80",X"32",X"22",X"84",X"32",X"2A",X"80",X"11",X"83",X"0D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"2A",X"80",X"A7",X"20",X"03",X"C3",X"E3",X"04",X"CD",X"F0",X"06",X"3A",
		X"28",X"80",X"3C",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",X"72",X"01",X"C3",
		X"E3",X"04",X"CD",X"00",X"10",X"3E",X"40",X"32",X"41",X"80",X"11",X"B3",X"0D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"3A",X"01",X"80",X"E6",X"07",X"C2",X"E6",X"04",X"21",X"41",X"80",X"35",X"28",
		X"03",X"C3",X"E6",X"04",X"3E",X"01",X"32",X"28",X"80",X"11",X"D6",X"04",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"C3",X"E3",X"04",X"CD",X"63",X"14",X"CD",X"27",X"14",X"C3",X"EF",X"12",X"D5",X"E5",
		X"5D",X"54",X"7D",X"CD",X"F2",X"0D",X"EB",X"7C",X"CD",X"F2",X"0D",X"19",X"CD",X"35",X"0E",X"E1",
		X"D1",X"C9",X"67",X"2E",X"00",X"CD",X"FB",X"0D",X"6C",X"67",X"C9",X"C5",X"D5",X"CD",X"12",X"0E",
		X"CB",X"79",X"28",X"06",X"47",X"7C",X"93",X"67",X"78",X"9A",X"CB",X"7A",X"28",X"01",X"91",X"D1",
		X"C1",X"C9",X"EB",X"4F",X"21",X"00",X"00",X"06",X"08",X"29",X"17",X"30",X"03",X"19",X"CE",X"00",
		X"10",X"F7",X"C9",X"C5",X"4F",X"AF",X"06",X"10",X"29",X"17",X"38",X"03",X"B9",X"38",X"02",X"91",
		X"23",X"10",X"F5",X"C1",X"C9",X"C5",X"D5",X"E5",X"06",X"08",X"11",X"40",X"00",X"7D",X"6C",X"62",
		X"A7",X"ED",X"52",X"30",X"01",X"19",X"3F",X"CB",X"12",X"87",X"ED",X"6A",X"87",X"ED",X"6A",X"10",
		X"EF",X"7A",X"E1",X"D1",X"C1",X"C9",X"C6",X"40",X"C5",X"E5",X"4F",X"CB",X"71",X"28",X"02",X"ED",
		X"44",X"E6",X"7F",X"21",X"71",X"0E",X"D7",X"7E",X"CB",X"79",X"28",X"02",X"ED",X"44",X"E1",X"C1",
		X"C9",X"00",X"03",X"06",X"09",X"0C",X"10",X"13",X"16",X"19",X"1C",X"1F",X"22",X"25",X"28",X"2B",
		X"2E",X"31",X"33",X"36",X"39",X"3C",X"3F",X"41",X"44",X"47",X"49",X"4C",X"4E",X"51",X"53",X"55",
		X"58",X"5A",X"5C",X"5E",X"60",X"62",X"64",X"66",X"68",X"6A",X"6B",X"6D",X"6F",X"70",X"71",X"73",
		X"74",X"75",X"76",X"78",X"79",X"7A",X"7A",X"7B",X"7C",X"7D",X"7D",X"7E",X"7E",X"7E",X"7F",X"7F",
		X"7F",X"7F",X"E5",X"CD",X"C4",X"0E",X"E1",X"CB",X"7D",X"28",X"03",X"2F",X"C6",X"81",X"CB",X"7C",
		X"C8",X"ED",X"44",X"C9",X"7C",X"DF",X"67",X"7D",X"DF",X"6F",X"BC",X"38",X"11",X"2E",X"00",X"CD",
		X"23",X"0E",X"29",X"29",X"29",X"29",X"29",X"7C",X"21",X"E7",X"0E",X"D7",X"7E",X"C9",X"7C",X"65",
		X"CD",X"CD",X"0E",X"2F",X"C6",X"41",X"C9",X"00",X"01",X"03",X"04",X"05",X"06",X"08",X"09",X"0A",
		X"0B",X"0C",X"0D",X"0F",X"10",X"11",X"12",X"13",X"14",X"15",X"16",X"17",X"18",X"19",X"19",X"1A",
		X"1B",X"1C",X"1D",X"1D",X"1E",X"1F",X"1F",X"20",X"CD",X"12",X"0F",X"CD",X"25",X"0F",X"CD",X"38",
		X"0F",X"C9",X"3A",X"85",X"80",X"A7",X"C8",X"21",X"80",X"80",X"01",X"07",X"68",X"CD",X"10",X"01",
		X"AF",X"32",X"85",X"80",X"C9",X"3A",X"95",X"80",X"A7",X"C8",X"21",X"90",X"80",X"01",X"07",X"68",
		X"CD",X"10",X"01",X"AF",X"32",X"95",X"80",X"C9",X"3A",X"A6",X"80",X"A7",X"C8",X"21",X"A0",X"80",
		X"01",X"08",X"68",X"CD",X"10",X"01",X"AF",X"32",X"A6",X"80",X"C9",X"E5",X"2A",X"08",X"80",X"7D",
		X"87",X"87",X"85",X"3C",X"6F",X"7C",X"E6",X"84",X"28",X"04",X"EE",X"84",X"20",X"01",X"37",X"7C",
		X"8F",X"67",X"85",X"22",X"08",X"80",X"E1",X"C9",X"3A",X"83",X"81",X"A7",X"C8",X"47",X"C5",X"3E",
		X"25",X"21",X"23",X"1B",X"E5",X"0E",X"C0",X"CD",X"5D",X"14",X"E1",X"C1",X"0E",X"B0",X"3E",X"2A",
		X"C3",X"5D",X"14",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"77",
		X"CD",X"0D",X"07",X"CD",X"2A",X"07",X"CD",X"AA",X"08",X"18",X"06",X"CD",X"0D",X"07",X"CD",X"47",
		X"07",X"CD",X"27",X"14",X"CD",X"EF",X"12",X"CD",X"63",X"14",X"21",X"15",X"16",X"11",X"B8",X"10",
		X"0E",X"C0",X"06",X"12",X"CD",X"1F",X"14",X"21",X"18",X"19",X"11",X"CA",X"10",X"06",X"03",X"CD",
		X"1F",X"14",X"26",X"14",X"11",X"12",X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"13",X"85",X"06",
		X"0A",X"CD",X"1F",X"14",X"21",X"1A",X"19",X"11",X"CD",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",
		X"14",X"11",X"22",X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"23",X"85",X"06",X"0A",X"CD",X"1F",
		X"14",X"21",X"1C",X"19",X"11",X"D0",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"32",
		X"85",X"CD",X"47",X"14",X"26",X"0B",X"11",X"33",X"85",X"06",X"0A",X"CD",X"1F",X"14",X"21",X"1E",
		X"19",X"11",X"D3",X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"42",X"85",X"CD",X"47",
		X"14",X"26",X"0B",X"11",X"43",X"85",X"06",X"0A",X"CD",X"1F",X"14",X"21",X"20",X"19",X"11",X"D6",
		X"10",X"06",X"03",X"CD",X"1F",X"14",X"26",X"14",X"11",X"52",X"85",X"CD",X"47",X"14",X"26",X"0B",
		X"11",X"53",X"85",X"06",X"0A",X"C3",X"1F",X"14",X"0B",X"3A",X"48",X"49",X"24",X"0F",X"3E",X"4B",
		X"3A",X"24",X"20",X"0A",X"1B",X"1B",X"12",X"18",X"1B",X"1C",X"01",X"48",X"49",X"02",X"43",X"39",
		X"03",X"47",X"39",X"04",X"49",X"3D",X"05",X"49",X"3D",X"21",X"F3",X"10",X"11",X"10",X"85",X"01",
		X"50",X"00",X"ED",X"B0",X"21",X"F0",X"10",X"11",X"24",X"80",X"01",X"03",X"00",X"ED",X"B0",X"C9",
		X"00",X"40",X"00",X"00",X"40",X"00",X"16",X"50",X"17",X"36",X"40",X"36",X"42",X"4A",X"47",X"36",
		X"00",X"00",X"00",X"00",X"35",X"00",X"0E",X"3E",X"47",X"47",X"4E",X"24",X"16",X"44",X"4A",X"50",
		X"00",X"00",X"00",X"00",X"30",X"00",X"0E",X"4B",X"3A",X"4F",X"44",X"44",X"24",X"0E",X"43",X"39",
		X"00",X"00",X"00",X"00",X"25",X"00",X"1C",X"50",X"18",X"40",X"36",X"42",X"44",X"49",X"44",X"24",
		X"00",X"00",X"00",X"00",X"20",X"00",X"1C",X"50",X"14",X"44",X"3F",X"3E",X"42",X"36",X"24",X"24",
		X"00",X"00",X"00",X"21",X"80",X"81",X"11",X"00",X"85",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"11",
		X"04",X"85",X"36",X"24",X"01",X"09",X"00",X"ED",X"B0",X"06",X"05",X"21",X"00",X"85",X"78",X"87",
		X"87",X"87",X"87",X"4F",X"C6",X"02",X"D7",X"11",X"02",X"85",X"1A",X"BE",X"38",X"23",X"20",X"0E",
		X"2D",X"1D",X"1A",X"BE",X"38",X"1B",X"20",X"06",X"2D",X"1D",X"1A",X"BE",X"38",X"13",X"21",X"00",
		X"85",X"79",X"D7",X"54",X"7D",X"C6",X"10",X"5F",X"C5",X"01",X"10",X"00",X"ED",X"B0",X"C1",X"10",
		X"CA",X"78",X"32",X"46",X"80",X"FE",X"05",X"CA",X"4E",X"06",X"21",X"10",X"85",X"07",X"07",X"07",
		X"07",X"D7",X"EB",X"21",X"00",X"85",X"01",X"10",X"00",X"ED",X"B0",X"CD",X"0B",X"10",X"CD",X"A1",
		X"12",X"26",X"19",X"3A",X"46",X"80",X"87",X"C6",X"18",X"6F",X"06",X"18",X"0E",X"B0",X"3E",X"1B",
		X"CD",X"5D",X"14",X"5D",X"16",X"0B",X"21",X"13",X"85",X"3A",X"46",X"80",X"87",X"87",X"87",X"87",
		X"85",X"6F",X"3E",X"0A",X"32",X"4D",X"80",X"3E",X"80",X"32",X"41",X"80",X"ED",X"53",X"50",X"80",
		X"22",X"52",X"80",X"F7",X"3A",X"00",X"A0",X"A7",X"20",X"78",X"3A",X"46",X"80",X"A7",X"28",X"02",
		X"3E",X"01",X"21",X"02",X"A0",X"D7",X"36",X"01",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",
		X"04",X"3A",X"21",X"80",X"D7",X"CB",X"66",X"28",X"41",X"CD",X"7F",X"12",X"2A",X"50",X"80",X"0E",
		X"C0",X"CD",X"4F",X"14",X"3A",X"01",X"80",X"4F",X"E6",X"07",X"C0",X"79",X"E6",X"1F",X"20",X"06",
		X"21",X"41",X"80",X"35",X"28",X"3C",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",X"04",X"3A",
		X"21",X"80",X"D7",X"7E",X"E6",X"0F",X"FE",X"02",X"28",X"38",X"FE",X"06",X"C0",X"2A",X"52",X"80",
		X"7E",X"3D",X"FE",X"09",X"20",X"02",X"3E",X"24",X"77",X"C9",X"CD",X"7F",X"12",X"77",X"23",X"22",
		X"52",X"80",X"2A",X"50",X"80",X"0E",X"C0",X"CD",X"4F",X"14",X"22",X"50",X"80",X"21",X"4D",X"80",
		X"35",X"C0",X"AF",X"32",X"02",X"A0",X"32",X"03",X"A0",X"32",X"16",X"A0",X"32",X"17",X"A0",X"C3",
		X"4E",X"06",X"2A",X"52",X"80",X"7E",X"3C",X"FE",X"25",X"20",X"02",X"3E",X"0A",X"77",X"C9",X"3A",
		X"20",X"80",X"A7",X"3A",X"16",X"80",X"28",X"0D",X"3A",X"21",X"80",X"A7",X"3A",X"16",X"80",X"28",
		X"04",X"0F",X"0F",X"0F",X"0F",X"0F",X"3E",X"00",X"38",X"02",X"3E",X"2C",X"2A",X"52",X"80",X"86",
		X"C9",X"21",X"09",X"15",X"11",X"CD",X"12",X"0E",X"C0",X"06",X"10",X"CD",X"1F",X"14",X"21",X"0C",
		X"16",X"11",X"DD",X"12",X"06",X"12",X"CD",X"1F",X"14",X"0E",X"B0",X"21",X"09",X"15",X"3E",X"1A",
		X"06",X"10",X"CD",X"5D",X"14",X"21",X"0C",X"16",X"06",X"12",X"C3",X"5D",X"14",X"0C",X"18",X"17",
		X"10",X"1B",X"0A",X"1D",X"1E",X"15",X"0A",X"1D",X"12",X"18",X"17",X"1C",X"2C",X"0E",X"17",X"1D",
		X"0E",X"1B",X"24",X"22",X"18",X"1E",X"1B",X"24",X"12",X"17",X"12",X"1D",X"12",X"0A",X"15",X"21",
		X"00",X"12",X"11",X"C3",X"3E",X"06",X"0A",X"0E",X"C0",X"CD",X"1F",X"14",X"21",X"00",X"12",X"06",
		X"0A",X"3E",X"1F",X"0E",X"B0",X"CD",X"5D",X"14",X"C9",X"01",X"99",X"03",X"2B",X"71",X"10",X"FC",
		X"C9",X"11",X"82",X"81",X"CD",X"1A",X"13",X"11",X"C2",X"81",X"21",X"26",X"80",X"06",X"03",X"1A",
		X"BE",X"D8",X"20",X"05",X"1B",X"2B",X"10",X"F7",X"C9",X"1A",X"77",X"1B",X"2B",X"10",X"FA",X"3A",
		X"21",X"80",X"3C",X"32",X"27",X"80",X"CD",X"63",X"14",X"C9",X"CD",X"27",X"14",X"CD",X"A9",X"13",
		X"3A",X"8C",X"81",X"A7",X"C0",X"ED",X"5B",X"89",X"81",X"2A",X"81",X"81",X"A7",X"ED",X"52",X"19",
		X"D8",X"3A",X"17",X"80",X"07",X"07",X"07",X"E6",X"03",X"28",X"02",X"3E",X"01",X"21",X"FB",X"13",
		X"CF",X"5E",X"23",X"56",X"EB",X"3A",X"17",X"80",X"2F",X"0F",X"0F",X"E6",X"07",X"CF",X"5E",X"23",
		X"56",X"2A",X"89",X"81",X"A7",X"ED",X"52",X"19",X"38",X"29",X"3A",X"17",X"80",X"2F",X"0F",X"0F",
		X"E6",X"07",X"FE",X"06",X"20",X"05",X"3E",X"01",X"32",X"8C",X"81",X"7D",X"83",X"27",X"6F",X"7C",
		X"8A",X"27",X"67",X"22",X"89",X"81",X"3A",X"83",X"81",X"3C",X"32",X"83",X"81",X"32",X"04",X"A0",
		X"C3",X"68",X"0F",X"ED",X"53",X"89",X"81",X"18",X"ED",X"21",X"81",X"81",X"7E",X"E6",X"F0",X"C8",
		X"0F",X"0F",X"0F",X"0F",X"4F",X"7E",X"E6",X"0F",X"C8",X"A1",X"C8",X"4F",X"2D",X"7E",X"E6",X"F0",
		X"C8",X"0F",X"0F",X"0F",X"0F",X"A1",X"C8",X"4F",X"7E",X"E6",X"0F",X"C8",X"A1",X"C8",X"3A",X"7E",
		X"79",X"FE",X"02",X"C0",X"21",X"CD",X"3E",X"11",X"E8",X"13",X"06",X"13",X"1A",X"07",X"2F",X"BE",
		X"C2",X"00",X"00",X"13",X"23",X"10",X"F5",X"C9",X"69",X"E8",X"EB",X"ED",X"7F",X"7B",X"FB",X"FE",
		X"ED",X"74",X"FA",X"F4",X"F9",X"F3",X"ED",X"75",X"71",X"79",X"D7",X"FF",X"13",X"0F",X"14",X"70",
		X"00",X"50",X"00",X"50",X"00",X"60",X"00",X"80",X"00",X"00",X"01",X"80",X"00",X"FF",X"FF",X"60",
		X"00",X"40",X"00",X"50",X"00",X"50",X"00",X"70",X"00",X"80",X"00",X"60",X"00",X"FF",X"FF",X"1A",
		X"CD",X"4F",X"14",X"13",X"10",X"F9",X"C9",X"0E",X"C0",X"21",X"01",X"1B",X"11",X"01",X"08",X"3A",
		X"21",X"80",X"A7",X"28",X"01",X"EB",X"D5",X"11",X"82",X"81",X"CD",X"47",X"14",X"E1",X"3A",X"22",
		X"80",X"A7",X"28",X"15",X"11",X"C2",X"81",X"06",X"03",X"3E",X"05",X"CD",X"6D",X"14",X"AF",X"E5",
		X"F5",X"CD",X"9B",X"14",X"F1",X"77",X"E1",X"25",X"C9",X"3E",X"24",X"06",X"07",X"CD",X"4F",X"14",
		X"10",X"FB",X"C9",X"0E",X"C0",X"21",X"01",X"11",X"11",X"26",X"80",X"18",X"DA",X"C5",X"47",X"1A",
		X"0F",X"0F",X"0F",X"0F",X"E6",X"0F",X"20",X"07",X"05",X"3E",X"24",X"F2",X"81",X"14",X"AF",X"06",
		X"00",X"CD",X"4F",X"14",X"1A",X"E6",X"0F",X"20",X"07",X"05",X"3E",X"24",X"F2",X"92",X"14",X"AF",
		X"06",X"00",X"CD",X"4F",X"14",X"78",X"C1",X"1B",X"10",X"D3",X"C9",X"3A",X"03",X"80",X"25",X"A7",
		X"3E",X"04",X"28",X"03",X"25",X"3E",X"18",X"85",X"E6",X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",
		X"67",X"E6",X"C0",X"B5",X"6F",X"7C",X"E6",X"07",X"81",X"67",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",
		X"C0",X"21",X"02",X"00",X"22",X"46",X"79",X"21",X"02",X"80",X"22",X"44",X"79",X"21",X"14",X"20",
		X"22",X"44",X"7C",X"21",X"50",X"01",X"22",X"46",X"7C",X"21",X"00",X"25",X"22",X"46",X"7A",X"21",
		X"00",X"0F",X"22",X"46",X"7B",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"CF",X"3A",X"28",X"80",X"A7",
		X"20",X"05",X"3E",X"01",X"32",X"0E",X"A0",X"CD",X"FE",X"15",X"CD",X"C1",X"15",X"CD",X"B8",X"16",
		X"CD",X"45",X"16",X"D0",X"AF",X"32",X"0E",X"A0",X"32",X"22",X"A0",X"3A",X"28",X"80",X"A7",X"20",
		X"0B",X"21",X"BA",X"15",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"3E",X"01",X"32",X"44",
		X"80",X"21",X"00",X"00",X"22",X"46",X"7D",X"21",X"C0",X"30",X"22",X"46",X"7C",X"F7",X"3A",X"2A",
		X"80",X"A7",X"20",X"87",X"3A",X"46",X"7D",X"3C",X"E6",X"07",X"32",X"46",X"7D",X"20",X"1F",X"3A",
		X"47",X"7D",X"3C",X"32",X"47",X"7D",X"FE",X"07",X"28",X"2A",X"FE",X"02",X"CC",X"A1",X"15",X"FE",
		X"04",X"CC",X"B1",X"15",X"FE",X"06",X"CC",X"A1",X"15",X"C6",X"30",X"32",X"47",X"7C",X"21",X"93",
		X"15",X"3A",X"47",X"7D",X"CF",X"3A",X"01",X"80",X"E6",X"0C",X"86",X"32",X"47",X"79",X"23",X"7E",
		X"32",X"46",X"7C",X"C9",X"3E",X"20",X"32",X"46",X"7D",X"AF",X"32",X"46",X"79",X"F7",X"21",X"46",
		X"7D",X"35",X"C0",X"21",X"8B",X"81",X"34",X"21",X"2A",X"80",X"36",X"01",X"AF",X"32",X"44",X"80",
		X"C3",X"BB",X"14",X"00",X"C0",X"00",X"C1",X"03",X"C4",X"03",X"C8",X"00",X"C2",X"00",X"C3",X"03",
		X"CC",X"21",X"47",X"7B",X"34",X"21",X"47",X"7A",X"35",X"F5",X"3E",X"2E",X"32",X"47",X"7C",X"F1",
		X"C9",X"21",X"47",X"7B",X"35",X"21",X"47",X"7A",X"34",X"C9",X"30",X"40",X"00",X"02",X"DF",X"10",
		X"10",X"2A",X"46",X"7A",X"3A",X"C6",X"7A",X"CF",X"11",X"00",X"12",X"A7",X"ED",X"52",X"19",X"30",
		X"01",X"EB",X"11",X"00",X"26",X"A7",X"ED",X"52",X"19",X"38",X"01",X"EB",X"22",X"46",X"7A",X"2A",
		X"46",X"7B",X"3A",X"C6",X"7B",X"CF",X"11",X"00",X"02",X"A7",X"ED",X"52",X"19",X"30",X"01",X"EB",
		X"11",X"00",X"1C",X"A7",X"ED",X"52",X"19",X"38",X"01",X"EB",X"22",X"46",X"7B",X"C9",X"3A",X"28",
		X"80",X"A7",X"20",X"1E",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",X"04",X"3A",X"21",X"80",
		X"D7",X"7E",X"E6",X"0F",X"21",X"33",X"16",X"CF",X"7E",X"32",X"C6",X"7A",X"23",X"7E",X"32",X"C6",
		X"7B",X"C9",X"3A",X"01",X"80",X"E6",X"0F",X"C0",X"CD",X"4B",X"0F",X"E6",X"0F",X"FE",X"09",X"30",
		X"F7",X"18",X"E1",X"F0",X"00",X"F0",X"F0",X"00",X"E8",X"10",X"F0",X"10",X"00",X"10",X"10",X"00",
		X"18",X"F0",X"10",X"00",X"00",X"ED",X"5B",X"46",X"82",X"3A",X"47",X"83",X"1F",X"CB",X"1A",X"FD",
		X"21",X"4E",X"79",X"06",X"19",X"CD",X"70",X"16",X"D8",X"FD",X"2C",X"FD",X"2C",X"10",X"F6",X"FD",
		X"21",X"20",X"79",X"06",X"10",X"CD",X"95",X"16",X"D8",X"FD",X"2C",X"FD",X"2C",X"10",X"F6",X"C9",
		X"3E",X"02",X"FD",X"BE",X"00",X"20",X"1C",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",
		X"96",X"D6",X"08",X"C6",X"10",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"04",
		X"C6",X"08",X"C9",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"F7",X"3E",X"09",X"FD",X"84",
		X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"1C",X"C6",X"28",X"D0",X"2C",X"24",X"7E",X"1F",X"25",
		X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"3A",X"42",X"79",X"FE",X"02",X"28",X"02",X"3E",
		X"01",X"C6",X"1F",X"4F",X"06",X"00",X"3A",X"01",X"80",X"E6",X"04",X"28",X"1B",X"ED",X"5B",X"44",
		X"82",X"3A",X"45",X"83",X"1F",X"CB",X"1A",X"FD",X"21",X"04",X"79",X"06",X"0E",X"CD",X"04",X"17",
		X"38",X"1C",X"FD",X"2C",X"FD",X"2C",X"10",X"F5",X"79",X"80",X"32",X"45",X"7C",X"3E",X"F4",X"2A",
		X"46",X"7A",X"84",X"67",X"22",X"44",X"7A",X"2A",X"46",X"7B",X"22",X"44",X"7B",X"C9",X"06",X"09",
		X"18",X"E6",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"F7",X"3E",X"09",X"FD",X"84",X"67",
		X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"0A",X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",
		X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"21",X"14",X"01",
		X"22",X"32",X"80",X"AF",X"32",X"30",X"80",X"21",X"A2",X"17",X"22",X"48",X"78",X"21",X"48",X"78",
		X"11",X"4A",X"78",X"01",X"04",X"00",X"ED",X"B0",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"D8",X"3A",
		X"44",X"80",X"A7",X"CC",X"72",X"17",X"DD",X"E5",X"DD",X"21",X"48",X"78",X"06",X"03",X"DD",X"5D",
		X"DD",X"54",X"CD",X"54",X"04",X"DD",X"2C",X"DD",X"2C",X"10",X"F3",X"DD",X"E1",X"AF",X"32",X"30",
		X"80",X"C9",X"3A",X"28",X"80",X"A7",X"20",X"23",X"3A",X"20",X"80",X"A7",X"21",X"19",X"80",X"28",
		X"04",X"3A",X"21",X"80",X"D7",X"CB",X"6E",X"21",X"33",X"80",X"28",X"03",X"36",X"01",X"C9",X"35",
		X"C0",X"3A",X"32",X"80",X"77",X"3E",X"01",X"32",X"30",X"80",X"C9",X"CD",X"4B",X"0F",X"E6",X"0F",
		X"18",X"E5",X"F7",X"EB",X"4C",X"11",X"30",X"80",X"1A",X"3D",X"C0",X"12",X"24",X"36",X"02",X"CB",
		X"FD",X"36",X"02",X"24",X"36",X"A0",X"3C",X"32",X"0B",X"A0",X"ED",X"5B",X"46",X"7A",X"CB",X"BD",
		X"73",X"2C",X"72",X"ED",X"5B",X"46",X"7B",X"24",X"72",X"2D",X"73",X"61",X"EB",X"F7",X"EB",X"C5",
		X"E5",X"CD",X"28",X"19",X"E1",X"C1",X"3A",X"01",X"80",X"F5",X"F5",X"E6",X"01",X"07",X"07",X"07",
		X"24",X"4C",X"2C",X"C6",X"80",X"77",X"F1",X"0F",X"E6",X"01",X"C6",X"23",X"24",X"24",X"24",X"77",
		X"F1",X"0F",X"0F",X"E6",X"01",X"C6",X"16",X"2D",X"77",X"61",X"7E",X"FE",X"03",X"28",X"0E",X"24",
		X"CD",X"4B",X"18",X"7A",X"FE",X"28",X"D8",X"25",X"2D",X"36",X"00",X"18",X"95",X"24",X"CB",X"FD",
		X"36",X"18",X"CB",X"BD",X"2C",X"24",X"24",X"36",X"23",X"2D",X"24",X"36",X"FF",X"F7",X"21",X"00",
		X"05",X"7C",X"DD",X"84",X"67",X"7D",X"DD",X"85",X"6F",X"34",X"7E",X"25",X"4C",X"25",X"25",X"25",
		X"FE",X"08",X"28",X"D5",X"F5",X"0F",X"E6",X"03",X"C6",X"18",X"61",X"77",X"F1",X"E6",X"01",X"07",
		X"07",X"07",X"25",X"25",X"25",X"2C",X"C6",X"80",X"77",X"2D",X"24",X"5E",X"2C",X"56",X"2D",X"CB",
		X"FD",X"EB",X"1A",X"CF",X"EB",X"CB",X"BD",X"73",X"2C",X"72",X"C9",X"CD",X"4B",X"0F",X"A7",X"C0",
		X"18",X"2A",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"44",X"80",X"A7",X"C0",X"3A",X"28",X"80",
		X"A7",X"20",X"E8",X"3A",X"20",X"80",X"A7",X"3A",X"16",X"80",X"28",X"0D",X"3A",X"21",X"80",X"A7",
		X"3A",X"16",X"80",X"28",X"04",X"0F",X"0F",X"0F",X"0F",X"0F",X"D8",X"F7",X"3A",X"40",X"79",X"FE",
		X"01",X"C0",X"F7",X"2A",X"46",X"7A",X"22",X"42",X"7A",X"3E",X"F4",X"84",X"67",X"22",X"40",X"7A",
		X"2A",X"46",X"7B",X"22",X"42",X"7B",X"22",X"40",X"7B",X"AF",X"32",X"C2",X"7A",X"32",X"42",X"7D",
		X"32",X"43",X"7D",X"3C",X"32",X"0C",X"A0",X"21",X"02",X"80",X"22",X"42",X"79",X"22",X"40",X"79",
		X"3E",X"1C",X"32",X"42",X"7C",X"21",X"14",X"22",X"22",X"40",X"7C",X"F7",X"21",X"42",X"7D",X"34",
		X"7E",X"E6",X"07",X"20",X"0C",X"2C",X"7E",X"FE",X"02",X"28",X"06",X"3C",X"77",X"25",X"2D",X"34",
		X"24",X"7E",X"0F",X"0F",X"E6",X"03",X"C6",X"25",X"32",X"43",X"7C",X"21",X"C2",X"7A",X"35",X"35",
		X"7E",X"2A",X"42",X"7A",X"CF",X"22",X"42",X"7A",X"2A",X"40",X"7A",X"3A",X"14",X"80",X"ED",X"44",
		X"CF",X"22",X"40",X"7A",X"CD",X"0B",X"19",X"D8",X"C3",X"62",X"18",X"2A",X"40",X"7A",X"ED",X"5B",
		X"42",X"7A",X"A7",X"ED",X"52",X"D8",X"AF",X"32",X"0C",X"A0",X"32",X"20",X"A0",X"CD",X"EE",X"19",
		X"AF",X"32",X"42",X"79",X"32",X"40",X"79",X"C9",X"3E",X"0A",X"DD",X"84",X"57",X"DD",X"5D",X"EB",
		X"5E",X"2C",X"56",X"24",X"7E",X"1F",X"CB",X"1A",X"FD",X"21",X"74",X"79",X"06",X"06",X"CD",X"A6",
		X"19",X"30",X"2F",X"FD",X"36",X"00",X"03",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"CB",X"FF",X"6F",
		X"36",X"00",X"3A",X"28",X"80",X"A7",X"20",X"1A",X"3E",X"03",X"FD",X"84",X"67",X"FD",X"7D",X"CB",
		X"FF",X"6F",X"7E",X"21",X"31",X"3D",X"D7",X"D5",X"C5",X"EB",X"E7",X"C1",X"D1",X"3E",X"01",X"32",
		X"05",X"A0",X"FD",X"2C",X"FD",X"2C",X"10",X"C6",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"CB",X"FF",
		X"6F",X"7E",X"CB",X"BD",X"77",X"FD",X"21",X"20",X"79",X"06",X"10",X"CD",X"CB",X"19",X"38",X"07",
		X"FD",X"2C",X"FD",X"2C",X"10",X"F5",X"C9",X"DD",X"7C",X"3C",X"67",X"DD",X"7D",X"6F",X"36",X"03",
		X"3E",X"01",X"32",X"0A",X"A0",X"C9",X"3E",X"02",X"FD",X"BE",X"00",X"20",X"1C",X"3E",X"09",X"FD",
		X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"10",X"C6",X"20",X"D0",X"2C",X"24",X"7E",X"1F",
		X"25",X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"A7",X"C9",X"3E",X"02",X"FD",X"BE",X"00",
		X"20",X"F7",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"18",X"C6",X"20",
		X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"08",X"C6",X"10",X"C9",X"ED",X"5B",
		X"40",X"82",X"3A",X"41",X"83",X"1F",X"CB",X"1A",X"FD",X"21",X"00",X"79",X"06",X"10",X"D5",X"CD",
		X"3D",X"1A",X"30",X"28",X"FD",X"36",X"00",X"03",X"3A",X"28",X"80",X"A7",X"20",X"1E",X"3E",X"03",
		X"FD",X"84",X"67",X"FD",X"7D",X"CB",X"FF",X"6F",X"7E",X"21",X"31",X"3D",X"D7",X"EB",X"C5",X"E7",
		X"21",X"36",X"1A",X"11",X"90",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C1",X"D1",X"FD",X"2C",X"FD",
		X"2C",X"10",X"CB",X"C9",X"A7",X"C9",X"40",X"40",X"40",X"01",X"FF",X"20",X"20",X"3E",X"02",X"FD",
		X"BE",X"00",X"20",X"F0",X"3E",X"09",X"FD",X"84",X"67",X"FD",X"7D",X"6F",X"7B",X"96",X"D6",X"0A",
		X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",X"25",X"7E",X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",
		X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"36",X"07",X"2D",X"36",
		X"17",X"CB",X"FD",X"36",X"0F",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",
		X"31",X"EB",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",
		X"2C",X"5D",X"36",X"03",X"2C",X"36",X"02",X"2C",X"36",X"00",X"24",X"36",X"01",X"24",X"16",X"7B",
		X"1A",X"3D",X"77",X"2D",X"1D",X"1A",X"77",X"24",X"36",X"17",X"2C",X"36",X"07",X"2D",X"CB",X"FD",
		X"36",X"1B",X"CB",X"BD",X"2D",X"2D",X"36",X"48",X"2C",X"2C",X"26",X"78",X"11",X"DD",X"1A",X"73",
		X"2C",X"72",X"11",X"CB",X"1A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",X"1C",
		X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",
		X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"16",X"32",X"EB",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",
		X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"2D",X"36",X"1F",X"CB",
		X"FD",X"36",X"15",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"11",X"26",X"7C",
		X"2C",X"3A",X"1C",X"80",X"77",X"EB",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"3A",
		X"88",X"81",X"D6",X"02",X"30",X"01",X"AF",X"32",X"88",X"81",X"C3",X"86",X"31",X"16",X"7E",X"DD",
		X"5D",X"3A",X"A3",X"81",X"12",X"16",X"79",X"18",X"10",X"16",X"7E",X"DD",X"5D",X"3A",X"B0",X"81",
		X"12",X"16",X"79",X"18",X"04",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",
		X"7C",X"2D",X"36",X"2C",X"CB",X"FD",X"36",X"1B",X"CB",X"BD",X"26",X"7E",X"CD",X"4B",X"0F",X"A6",
		X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",
		X"7A",X"2C",X"3A",X"B1",X"81",X"BE",X"38",X"64",X"2D",X"26",X"7D",X"3A",X"01",X"80",X"E6",X"07",
		X"20",X"37",X"35",X"20",X"34",X"11",X"8E",X"1B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",X"7D",X"34",X"7E",X"FE",X"0C",X"20",
		X"06",X"E5",X"CD",X"87",X"32",X"E1",X"7E",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1A",X"EB",
		X"21",X"F9",X"1B",X"D7",X"15",X"7E",X"12",X"14",X"EB",X"2C",X"25",X"3A",X"1C",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"24",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",
		X"77",X"11",X"64",X"1B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"18",X"DD",X"11",X"E5",X"1B",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",
		X"EB",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"2D",X"2E",X"2F",X"2E",X"2D",X"2C",
		X"16",X"7E",X"DD",X"5D",X"3A",X"A0",X"81",X"12",X"16",X"79",X"18",X"10",X"16",X"7E",X"DD",X"5D",
		X"3A",X"B0",X"81",X"12",X"16",X"79",X"18",X"04",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7C",X"2D",X"36",X"27",X"CB",X"FD",X"36",X"30",X"CB",X"BD",X"26",X"7E",X"CD",
		X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"86",X"31",X"26",X"7D",X"16",X"7A",X"5D",X"1C",X"1A",X"4F",X"3A",X"B1",X"81",X"B9",X"D4",X"71",
		X"32",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",
		X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"5D",X"36",X"03",X"2C",X"36",X"02",X"2C",
		X"36",X"00",X"24",X"36",X"01",X"24",X"16",X"7B",X"1A",X"3D",X"77",X"2D",X"1D",X"1A",X"77",X"24",
		X"36",X"27",X"CB",X"FD",X"36",X"36",X"CB",X"BD",X"2D",X"2D",X"36",X"44",X"2C",X"2C",X"26",X"7E",
		X"3A",X"A0",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",X"78",X"11",X"BE",X"1C",
		X"73",X"2C",X"72",X"11",X"AC",X"1C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",
		X"1C",X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"16",X"32",X"26",X"7D",X"CD",X"71",X"32",X"25",X"2C",
		X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"C5",X"16",
		X"78",X"DD",X"5D",X"D5",X"21",X"47",X"1D",X"01",X"0A",X"00",X"ED",X"B0",X"D1",X"14",X"D5",X"6B",
		X"62",X"36",X"02",X"2C",X"36",X"00",X"2C",X"EB",X"01",X"08",X"00",X"ED",X"B0",X"D1",X"D5",X"CB",
		X"FB",X"7B",X"C6",X"08",X"EB",X"E5",X"77",X"2C",X"36",X"7C",X"2C",X"EB",X"E1",X"01",X"06",X"00",
		X"ED",X"B0",X"D1",X"14",X"D5",X"21",X"51",X"1D",X"01",X"0A",X"00",X"ED",X"B0",X"D1",X"14",X"EB",
		X"4E",X"2C",X"46",X"2C",X"3E",X"80",X"81",X"F5",X"77",X"2C",X"70",X"F1",X"30",X"01",X"34",X"34",
		X"2C",X"79",X"D6",X"80",X"F5",X"77",X"2C",X"70",X"F1",X"30",X"01",X"35",X"35",X"2C",X"71",X"2C",
		X"70",X"2C",X"71",X"2C",X"70",X"C1",X"C9",X"9E",X"1D",X"9E",X"1D",X"9E",X"1D",X"9E",X"1D",X"5B",
		X"1D",X"00",X"00",X"80",X"01",X"80",X"01",X"00",X"03",X"80",X"01",X"16",X"7C",X"DD",X"5D",X"EB",
		X"36",X"3A",X"CB",X"FD",X"36",X"36",X"11",X"6F",X"1D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",
		X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"11",X"26",X"7C",X"2C",X"3A",X"1C",X"80",X"77",
		X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"54",X"5D",X"3E",X"03",X"2D",X"2D",
		X"77",X"2D",X"2D",X"77",X"2D",X"2D",X"77",X"2D",X"2D",X"77",X"EB",X"C3",X"86",X"31",X"16",X"7C",
		X"DD",X"5D",X"EB",X"26",X"7C",X"36",X"2C",X"CB",X"FD",X"36",X"1B",X"CB",X"BD",X"26",X"7E",X"3A",
		X"A5",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",
		X"7E",X"FE",X"03",X"28",X"59",X"26",X"7A",X"2C",X"3A",X"B1",X"81",X"BE",X"38",X"70",X"2D",X"26",
		X"7D",X"3A",X"01",X"80",X"E6",X"07",X"20",X"36",X"35",X"20",X"33",X"11",X"E4",X"1D",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"30",X"26",X"7D",
		X"34",X"7E",X"FE",X"0C",X"20",X"06",X"E5",X"CD",X"87",X"32",X"E1",X"7E",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"27",X"EB",X"21",X"5A",X"1E",X"D7",X"15",X"7E",X"12",X"14",X"EB",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"E5",X"CB",
		X"FD",X"5E",X"2C",X"56",X"EB",X"36",X"24",X"E1",X"C3",X"86",X"31",X"24",X"CD",X"4B",X"0F",X"A6",
		X"3C",X"25",X"77",X"11",X"BB",X"1D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"18",X"D0",X"11",X"47",
		X"1E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",
		X"CD",X"EB",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"2D",X"2E",X"2F",X"2E",X"2D",
		X"2C",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"2D",X"26",X"7C",X"36",X"00",
		X"CB",X"FD",X"36",X"36",X"F7",X"16",X"79",X"DD",X"5D",X"1A",X"FE",X"03",X"28",X"07",X"14",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"EB",X"26",X"7D",X"36",X"FF",X"11",X"93",X"1E",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"0F",X"0F",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"24",X"FE",X"04",X"20",X"08",X"26",X"79",X"2C",X"36",X"03",X"2D",X"26",X"7D",
		X"25",X"EB",X"21",X"F1",X"1E",X"D7",X"7E",X"EB",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",
		X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"79",X"36",X"02",X"11",X"D5",X"1E",X"DD",
		X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",
		X"EB",X"1C",X"16",X"7C",X"3A",X"1C",X"80",X"12",X"1D",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",
		X"30",X"A8",X"A9",X"AA",X"AB",X"AE",X"B2",X"B6",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"26",
		X"7C",X"36",X"15",X"2C",X"36",X"26",X"2D",X"CB",X"FD",X"36",X"21",X"F7",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"24",X"2C",X"3A",X"47",X"7A",X"BE",X"CB",X"FD",X"3E",X"00",X"38",X"35",X"28",
		X"02",X"3C",X"3C",X"77",X"CB",X"BD",X"24",X"3A",X"47",X"7B",X"BE",X"3E",X"00",X"38",X"29",X"28",
		X"02",X"3C",X"3C",X"2D",X"CB",X"FD",X"86",X"77",X"25",X"2C",X"7E",X"2D",X"86",X"77",X"CB",X"BD",
		X"26",X"79",X"2C",X"3A",X"01",X"80",X"E6",X"0C",X"C6",X"80",X"77",X"2D",X"24",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"3D",X"3D",X"18",X"CB",X"3D",X"3D",X"18",X"D7",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7B",X"CD",X"98",X"33",X"24",X"2D",X"36",X"00",X"CB",
		X"FD",X"36",X"30",X"11",X"7C",X"1F",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"1A",X"FE",X"03",X"28",X"08",X"16",X"7A",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"EB",X"2C",X"36",
		X"80",X"26",X"7C",X"36",X"0E",X"2D",X"36",X"1F",X"F7",X"CD",X"D6",X"1F",X"38",X"0A",X"16",X"7A",
		X"DD",X"5D",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"3A",X"16",X"80",X"CB",X"4F",X"20",X"08",X"11",
		X"70",X"3D",X"C5",X"E7",X"C1",X"18",X"0C",X"3A",X"83",X"81",X"3C",X"32",X"83",X"81",X"C5",X"CD",
		X"68",X"0F",X"C1",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"00",X"26",X"7F",X"36",X"00",X"3E",X"01",
		X"32",X"0D",X"A0",X"C3",X"79",X"30",X"16",X"82",X"DD",X"5D",X"EB",X"ED",X"5B",X"46",X"82",X"3A",
		X"47",X"83",X"1F",X"CB",X"1A",X"7B",X"96",X"D6",X"0A",X"C6",X"14",X"D0",X"2C",X"24",X"7E",X"1F",
		X"25",X"7E",X"1F",X"92",X"D6",X"05",X"C6",X"0A",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FB",
		X"CD",X"A7",X"20",X"F7",X"CD",X"CB",X"20",X"38",X"1A",X"24",X"3A",X"1C",X"80",X"77",X"2D",X"26",
		X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"A7",X"20",X"F7",X"CD",X"CB",X"20",X"38",
		X"71",X"18",X"E6",X"D6",X"02",X"38",X"38",X"11",X"30",X"20",X"DD",X"73",X"00",X"DD",X"72",X"01",
		X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",
		X"E6",X"07",X"EB",X"21",X"9F",X"20",X"D7",X"EB",X"25",X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",
		X"2D",X"25",X"CB",X"FD",X"35",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"11",
		X"68",X"20",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",
		X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"E6",X"07",X"C6",X"08",X"25",X"77",X"2C",X"3A",
		X"1C",X"80",X"77",X"2D",X"25",X"CB",X"FD",X"34",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",
		X"79",X"30",X"E5",X"F5",X"CD",X"87",X"32",X"F1",X"E1",X"D6",X"02",X"38",X"C2",X"18",X"88",X"0F",
		X"0E",X"0D",X"0C",X"0B",X"0A",X"09",X"08",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"06",X"CB",X"BD",X"36",X"08",X"24",X"36",X"00",X"C9",X"16",X"79",X"DD",X"5D",X"EB",
		X"7E",X"FE",X"03",X"CA",X"E2",X"20",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"02",X"C6",
		X"04",X"C9",X"33",X"33",X"C3",X"1F",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"8B",X"33",X"EB",X"15",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"09",X"CB",X"BD",X"36",X"10",X"24",X"CD",X"4B",X"0F",X"E6",X"3F",X"C6",X"40",X"77",
		X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"35",X"28",
		X"10",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"E5",X"CD",X"87",X"32",X"E1",X"11",X"3F",X"21",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",
		X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"0F",
		X"E6",X"0F",X"FE",X"07",X"28",X"13",X"C6",X"10",X"25",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"2C",X"26",X"7A",X"EB",X"1A",X"4F",X"3A",
		X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",X"CB",
		X"FB",X"1D",X"21",X"B3",X"3D",X"C6",X"80",X"CD",X"7E",X"33",X"EB",X"CB",X"BD",X"26",X"78",X"11",
		X"95",X"21",X"73",X"2C",X"72",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",
		X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"24",X"36",X"28",X"24",X"CD",
		X"98",X"33",X"18",X"0F",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7B",
		X"CD",X"8B",X"33",X"25",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",X"7C",X"36",X"0F",
		X"CB",X"BD",X"26",X"7E",X"3A",X"A4",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"F7",
		X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"3A",X"01",X"80",
		X"E6",X"07",X"20",X"1A",X"35",X"20",X"17",X"E5",X"CD",X"4B",X"0F",X"24",X"A6",X"3C",X"25",X"77",
		X"26",X"7A",X"2C",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"CD",X"87",X"32",X"E1",X"25",X"3A",
		X"01",X"80",X"E6",X"03",X"C6",X"28",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"00",
		X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"33",X"3E",X"CD",X"65",X"33",X"EB",X"26",X"7C",
		X"36",X"0C",X"CB",X"BD",X"26",X"7E",X"3A",X"A4",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",
		X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"3A",
		X"01",X"80",X"E6",X"07",X"20",X"1E",X"35",X"20",X"1B",X"E5",X"CD",X"4B",X"0F",X"24",X"A6",X"3C",
		X"25",X"77",X"26",X"7B",X"CB",X"FD",X"EB",X"CD",X"4B",X"0F",X"21",X"33",X"3E",X"CD",X"7E",X"33",
		X"CD",X"87",X"32",X"E1",X"25",X"3A",X"01",X"80",X"E6",X"03",X"C6",X"28",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"68",X"23",X"F7",
		X"CD",X"8C",X"23",X"38",X"0F",X"24",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"D6",X"06",X"38",X"56",X"11",X"D1",X"22",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"34",X"7E",
		X"0F",X"E6",X"07",X"FE",X"06",X"20",X"02",X"AF",X"77",X"EB",X"21",X"5C",X"23",X"D7",X"EB",X"25",
		X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"25",X"CB",X"FD",X"35",X"CB",X"BD",X"25",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"68",X"23",X"F7",X"CD",X"8C",X"23",X"38",X"02",X"18",
		X"A4",X"E5",X"F5",X"CD",X"87",X"32",X"F1",X"E1",X"D6",X"06",X"38",X"02",X"18",X"AA",X"11",X"27",
		X"23",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"34",X"7E",X"0F",X"E6",X"07",X"FE",X"06",X"20",X"02",X"AF",X"77",X"EB",
		X"21",X"62",X"23",X"D7",X"EB",X"25",X"1A",X"77",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"25",X"CB",
		X"FD",X"34",X"CB",X"BD",X"25",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"A0",X"A1",X"A2",X"A3",
		X"A4",X"A5",X"A5",X"A4",X"A3",X"A2",X"A1",X"A0",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"B3",X"3D",X"CD",X"65",X"33",X"EB",
		X"26",X"7C",X"36",X"12",X"CB",X"BD",X"36",X"A0",X"24",X"36",X"00",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"A3",X"23",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"06",
		X"C6",X"0C",X"C9",X"33",X"33",X"C3",X"1F",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",
		X"36",X"00",X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"EB",
		X"26",X"7C",X"36",X"1B",X"CB",X"BD",X"36",X"20",X"24",X"CD",X"4B",X"0F",X"E6",X"3F",X"C6",X"30",
		X"77",X"24",X"3A",X"A1",X"81",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"2C",X"36",X"00",X"26",X"7B",X"3A",X"47",X"7B",X"BE",
		X"3E",X"01",X"38",X"02",X"3E",X"FF",X"CB",X"FD",X"77",X"CB",X"BD",X"2D",X"26",X"7D",X"36",X"01",
		X"CD",X"71",X"32",X"11",X"1C",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"34",X"7E",X"0F",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1D",X"C6",X"20",X"2D",X"25",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",X"EB",X"CD",
		X"91",X"30",X"C3",X"79",X"30",X"11",X"5E",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",
		X"00",X"26",X"7B",X"CD",X"98",X"33",X"EB",X"15",X"21",X"B3",X"3D",X"CD",X"65",X"33",X"EB",X"26",
		X"7C",X"36",X"27",X"CB",X"BD",X"36",X"01",X"26",X"7E",X"3A",X"A2",X"81",X"77",X"CD",X"4B",X"0F",
		X"A6",X"25",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",
		X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"D6",X"04",X"C6",X"08",X"38",X"16",X"2D",X"26",X"7D",X"CD",
		X"71",X"32",X"25",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",
		X"79",X"30",X"D6",X"04",X"3E",X"02",X"38",X"02",X"3E",X"FE",X"CB",X"FD",X"77",X"CB",X"BD",X"26",
		X"7D",X"36",X"FF",X"11",X"FC",X"24",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",
		X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"34",X"7E",X"0F",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"1D",X"C6",X"01",X"2D",X"25",X"77",X"2C",X"3A",X"1C",
		X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",X"EB",X"CD",
		X"91",X"30",X"C3",X"79",X"30",X"11",X"3E",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",
		X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",X"CD",X"71",X"32",X"2C",X"25",
		X"3A",X"1C",X"80",X"77",X"CB",X"FD",X"25",X"7E",X"2D",X"86",X"77",X"25",X"35",X"35",X"CB",X"BD",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"0F",X"25",X"36",X"00",X"25",
		X"36",X"10",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",X"4B",
		X"0F",X"E6",X"FF",X"3C",X"77",X"25",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",X"02",
		X"11",X"99",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",
		X"03",X"CA",X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",
		X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"36",X"FF",X"26",X"79",X"36",X"03",X"CD",
		X"87",X"32",X"11",X"CB",X"25",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"A8",X"27",X"D2",X"9D",
		X"27",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"15",X"25",X"36",X"00",X"25",
		X"36",X"10",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7C",
		X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",X"02",X"11",X"03",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7B",
		X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"38",X"9B",X"25",X"2C",
		X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",
		X"28",X"36",X"12",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"CD",
		X"4B",X"0F",X"E6",X"3F",X"3C",X"77",X"25",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",
		X"02",X"2C",X"24",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"11",X"63",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7D",
		X"35",X"CA",X"B9",X"25",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",
		X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"1B",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"26",X"7C",X"36",X"11",X"2C",X"26",X"79",X"36",X"80",X"2D",X"36",
		X"02",X"2C",X"24",X"EB",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"11",X"B3",X"26",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",X"31",X"26",X"7B",
		X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"DA",X"B9",X"25",X"25",
		X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",
		X"26",X"28",X"36",X"24",X"F7",X"CD",X"E7",X"27",X"30",X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",
		X"CD",X"4B",X"0F",X"E6",X"3F",X"3C",X"77",X"25",X"36",X"12",X"2C",X"26",X"7A",X"EB",X"21",X"F3",
		X"3D",X"CD",X"65",X"33",X"EB",X"CB",X"BD",X"25",X"36",X"02",X"2C",X"36",X"80",X"11",X"16",X"27",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",
		X"31",X"26",X"7D",X"35",X"28",X"6B",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"CD",X"26",X"28",X"36",X"33",X"F7",X"CD",X"E7",X"27",X"30",
		X"06",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"25",X"36",X"12",X"2C",X"26",X"7A",X"EB",X"21",X"F3",
		X"3D",X"CD",X"65",X"33",X"EB",X"CB",X"BD",X"25",X"36",X"02",X"2C",X"36",X"80",X"11",X"66",X"27",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"1F",
		X"31",X"26",X"7B",X"2C",X"3A",X"47",X"7B",X"96",X"2D",X"26",X"7D",X"D6",X"04",X"C6",X"08",X"38",
		X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"36",X"FF",X"26",X"79",X"36",X"03",X"CD",X"D9",X"32",X"C3",X"C2",X"25",X"26",X"7F",X"36",
		X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",
		X"10",X"20",X"09",X"2C",X"26",X"7A",X"35",X"24",X"34",X"2D",X"26",X"7D",X"4F",X"0F",X"0F",X"E6",
		X"07",X"FE",X"05",X"D0",X"EB",X"21",X"DB",X"27",X"CF",X"15",X"7E",X"12",X"23",X"1C",X"16",X"79",
		X"79",X"07",X"07",X"E6",X"0C",X"86",X"12",X"1D",X"14",X"37",X"C9",X"04",X"80",X"05",X"80",X"06",
		X"80",X"07",X"80",X"08",X"83",X"0C",X"83",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",X"08",
		X"20",X"09",X"2C",X"26",X"7A",X"34",X"24",X"35",X"2D",X"26",X"7D",X"4F",X"0F",X"0F",X"E6",X"07",
		X"FE",X"05",X"D0",X"EB",X"21",X"1A",X"28",X"CF",X"15",X"7E",X"12",X"23",X"1C",X"16",X"79",X"79",
		X"07",X"07",X"E6",X"0C",X"86",X"12",X"1D",X"14",X"37",X"C9",X"0C",X"83",X"08",X"83",X"07",X"80",
		X"06",X"80",X"05",X"80",X"04",X"80",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"24",X"CD",
		X"4B",X"0F",X"E6",X"0F",X"C6",X"05",X"77",X"24",X"CD",X"8B",X"33",X"34",X"24",X"36",X"24",X"2D",
		X"24",X"36",X"FF",X"25",X"CB",X"FD",X"3E",X"01",X"32",X"09",X"A0",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"80",X"26",X"7B",X"CD",X"8B",X"33",X"24",X"2D",X"36",X"13",X"CB",
		X"FD",X"36",X"30",X"26",X"7A",X"36",X"30",X"24",X"36",X"00",X"CB",X"BD",X"26",X"7D",X"CD",X"4B",
		X"0F",X"E6",X"1F",X"C6",X"20",X"77",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"1F",X"31",X"26",X"7D",X"35",X"28",X"10",X"25",X"2C",X"3A",X"43",X"80",X"77",X"2D",X"26",X"7A",
		X"EB",X"CD",X"91",X"30",X"C3",X"79",X"30",X"E5",X"CD",X"0A",X"33",X"3E",X"01",X"32",X"06",X"A0",
		X"C5",X"21",X"B9",X"28",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C1",X"E1",X"26",X"7F",
		X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"30",X"80",X"80",X"01",X"FF",X"10",X"10",
		X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"EB",X"21",X"D9",X"28",X"3A",X"01",X"80",X"0F",X"E6",
		X"03",X"D7",X"7E",X"12",X"16",X"7A",X"C3",X"FC",X"30",X"32",X"33",X"30",X"31",X"16",X"79",X"DD",
		X"5D",X"EB",X"36",X"03",X"2C",X"36",X"00",X"26",X"7B",X"36",X"1E",X"F7",X"16",X"7A",X"DD",X"5D",
		X"1C",X"1A",X"4F",X"3A",X"47",X"7A",X"D6",X"02",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",
		X"D6",X"02",X"91",X"67",X"CD",X"B2",X"0E",X"CB",X"FB",X"1D",X"21",X"73",X"3D",X"CD",X"7E",X"33",
		X"CB",X"BB",X"1C",X"EB",X"3A",X"47",X"7A",X"D6",X"02",X"BE",X"20",X"A4",X"24",X"3A",X"47",X"7B",
		X"D6",X"02",X"BE",X"20",X"9B",X"11",X"2E",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",
		X"80",X"A7",X"20",X"06",X"3A",X"2E",X"80",X"A7",X"20",X"16",X"CD",X"F7",X"29",X"14",X"21",X"D9",
		X"28",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"C9",
		X"11",X"59",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"F7",X"29",X"3A",X"01",X"80",X"0F",
		X"0F",X"E6",X"07",X"FE",X"07",X"28",X"14",X"21",X"74",X"29",X"D7",X"14",X"7E",X"12",X"1C",X"3A",
		X"1C",X"80",X"12",X"C9",X"32",X"32",X"32",X"32",X"34",X"35",X"36",X"16",X"7D",X"EB",X"36",X"E0",
		X"11",X"89",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"28",
		X"20",X"EB",X"2A",X"46",X"7B",X"1A",X"D5",X"EF",X"D1",X"16",X"7B",X"EB",X"73",X"2C",X"72",X"ED",
		X"5B",X"46",X"7A",X"25",X"15",X"15",X"72",X"2D",X"73",X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",
		X"C9",X"26",X"7A",X"ED",X"5B",X"46",X"7A",X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",
		X"7B",X"72",X"2D",X"73",X"CB",X"FD",X"36",X"00",X"25",X"36",X"A0",X"3E",X"01",X"32",X"08",X"A0",
		X"11",X"D9",X"29",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7C",X"DD",X"5D",X"21",X"D9",X"28",
		X"3A",X"01",X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"1D",X"16",
		X"7A",X"CD",X"91",X"30",X"C3",X"79",X"30",X"16",X"7A",X"DD",X"5D",X"EB",X"ED",X"5B",X"46",X"7A",
		X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",X"7B",X"15",X"15",X"72",X"2D",X"73",X"EB",
		X"C9",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"2D",X"EB",X"21",X"2A",X"2A",X"3A",X"01",X"80",X"0F",
		X"E6",X"03",X"D7",X"7E",X"12",X"16",X"7A",X"C3",X"FC",X"30",X"32",X"31",X"30",X"33",X"16",X"79",
		X"DD",X"5D",X"EB",X"36",X"03",X"2C",X"36",X"00",X"F7",X"16",X"7A",X"DD",X"5D",X"1C",X"1A",X"4F",
		X"3A",X"47",X"7A",X"D6",X"02",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"C6",X"02",X"91",
		X"67",X"CD",X"B2",X"0E",X"CB",X"FB",X"1D",X"21",X"73",X"3D",X"CD",X"7E",X"33",X"CB",X"BB",X"1C",
		X"EB",X"3A",X"47",X"7A",X"D6",X"02",X"BE",X"20",X"A8",X"24",X"3A",X"47",X"7B",X"C6",X"02",X"BE",
		X"20",X"9F",X"11",X"7B",X"2A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"01",X"80",X"A7",X"20",
		X"06",X"3A",X"2E",X"80",X"A7",X"20",X"16",X"CD",X"09",X"2B",X"14",X"21",X"2A",X"2A",X"3A",X"01",
		X"80",X"0F",X"E6",X"03",X"D7",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",X"C9",X"11",X"A6",X"2A",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"09",X"2B",X"3A",X"01",X"80",X"0F",X"0F",X"E6",X"07",
		X"FE",X"07",X"28",X"14",X"21",X"C1",X"2A",X"D7",X"14",X"7E",X"12",X"1C",X"3A",X"1C",X"80",X"12",
		X"C9",X"32",X"32",X"32",X"32",X"37",X"38",X"39",X"16",X"7D",X"EB",X"36",X"20",X"11",X"D6",X"2A",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"35",X"28",X"20",X"EB",X"2A",
		X"46",X"7B",X"1A",X"D5",X"EF",X"D1",X"16",X"7B",X"EB",X"73",X"2C",X"72",X"ED",X"5B",X"46",X"7A",
		X"15",X"15",X"25",X"72",X"2D",X"73",X"2C",X"26",X"7C",X"3A",X"1C",X"80",X"77",X"C9",X"26",X"7F",
		X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",X"30",X"16",X"7A",X"DD",X"5D",X"EB",X"ED",X"5B",
		X"46",X"7A",X"15",X"15",X"73",X"2C",X"72",X"24",X"ED",X"5B",X"46",X"7B",X"14",X"14",X"72",X"2D",
		X"73",X"EB",X"C9",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"2C",X"36",X"82",X"24",X"2D",X"CB",
		X"FD",X"36",X"10",X"CB",X"BD",X"24",X"2C",X"CD",X"8B",X"33",X"34",X"F7",X"16",X"7A",X"DD",X"5D",
		X"EB",X"E5",X"7E",X"2C",X"17",X"7E",X"17",X"E6",X"07",X"EB",X"21",X"5D",X"2B",X"CF",X"7E",X"16",
		X"7C",X"12",X"23",X"7E",X"1D",X"12",X"D1",X"CD",X"D4",X"30",X"C3",X"79",X"30",X"2B",X"20",X"2C",
		X"21",X"2B",X"24",X"2C",X"25",X"2B",X"28",X"2C",X"29",X"2B",X"2C",X"2C",X"2D",X"16",X"7A",X"DD",
		X"5D",X"1C",X"21",X"F3",X"3D",X"CD",X"65",X"33",X"F7",X"16",X"7A",X"DD",X"5D",X"CD",X"91",X"30",
		X"C3",X"79",X"30",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"15",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",
		X"45",X"2E",X"26",X"7C",X"18",X"3F",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"1E",X"F7",X"CD",X"45",
		X"2E",X"CD",X"65",X"2E",X"18",X"2F",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"24",X"CB",X"BD",X"36",
		X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"BB",X"2E",X"38",X"04",X"26",X"7C",X"18",X"18",X"26",X"7A",
		X"CB",X"FD",X"36",X"0E",X"11",X"CD",X"2B",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",
		X"CD",X"65",X"2E",X"18",X"00",X"2C",X"3A",X"1C",X"80",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"D4",
		X"30",X"C3",X"79",X"30",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"2A",X"CB",X"BD",X"36",X"4C",X"F7",
		X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"04",X"26",X"7C",X"18",X"DA",X"26",X"7A",X"CB",X"FD",
		X"36",X"0E",X"11",X"0B",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",
		X"35",X"28",X"05",X"CD",X"65",X"2E",X"18",X"BD",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"27",
		X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7C",X"18",X"A7",X"0E",X"0E",
		X"CD",X"8C",X"2E",X"36",X"30",X"F7",X"CD",X"45",X"2E",X"CD",X"BB",X"2E",X"38",X"06",X"2D",X"CD",
		X"65",X"2E",X"18",X"91",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"53",X"2C",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"04",X"25",X"C3",X"D5",X"2B",X"26",
		X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"6E",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",
		X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"33",X"CB",X"BD",
		X"36",X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"05",X"26",X"7C",X"C3",X"D6",X"2B",
		X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"9F",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",
		X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",
		X"FD",X"36",X"08",X"11",X"BC",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",
		X"7C",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"36",X"F7",X"CD",X"45",X"2E",X"CD",
		X"BB",X"2E",X"38",X"07",X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",
		X"16",X"11",X"EA",X"2C",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",
		X"28",X"06",X"CD",X"81",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"07",
		X"2D",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",
		X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"39",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"07",
		X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"36",X"2D",
		X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",
		X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"53",X"2D",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"CD",X"45",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",
		X"2E",X"36",X"3F",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",X"45",X"2E",X"CD",X"A0",X"2E",X"38",X"05",
		X"26",X"7C",X"C3",X"D6",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"16",X"11",X"84",X"2D",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"CD",X"45",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"81",X"2E",X"C3",
		X"D5",X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"08",X"11",X"68",X"2D",X"DD",X"73",X"00",X"DD",X"72",
		X"01",X"18",X"C5",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"15",X"CB",X"BD",X"36",X"4C",X"F7",X"CD",
		X"55",X"2E",X"26",X"7C",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"1E",X"F7",X"CD",
		X"55",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"08",X"CD",X"8C",X"2E",X"36",X"24",X"CB",
		X"BD",X"36",X"4C",X"F7",X"CD",X"55",X"2E",X"CD",X"BB",X"2E",X"38",X"05",X"26",X"7C",X"C3",X"D6",
		X"2B",X"26",X"7A",X"CB",X"FD",X"36",X"0E",X"11",X"F0",X"2D",X"DD",X"73",X"00",X"DD",X"72",X"01",
		X"CD",X"55",X"2E",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",X"0E",X"0E",X"CD",X"8C",X"2E",X"36",X"39",
		X"F7",X"CD",X"55",X"2E",X"CD",X"A0",X"2E",X"38",X"07",X"2D",X"CD",X"65",X"2E",X"C3",X"D5",X"2B",
		X"26",X"7A",X"CB",X"FD",X"36",X"02",X"11",X"1F",X"2E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",
		X"55",X"2E",X"26",X"7D",X"35",X"28",X"06",X"CD",X"71",X"2E",X"C3",X"D5",X"2B",X"26",X"7A",X"CB",
		X"FD",X"36",X"0E",X"11",X"3C",X"2E",X"DD",X"73",X"00",X"DD",X"72",X"01",X"CD",X"55",X"2E",X"CD",
		X"65",X"2E",X"C3",X"D5",X"2B",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"01",X"C9",
		X"33",X"33",X"C3",X"86",X"31",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"28",X"01",X"C9",
		X"33",X"33",X"C3",X"16",X"32",X"26",X"7C",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"C6",X"4C",X"77",
		X"C9",X"26",X"7C",X"3A",X"01",X"80",X"0F",X"E6",X"03",X"ED",X"44",X"E6",X"03",X"C6",X"4C",X"77",
		X"C9",X"26",X"7C",X"3A",X"01",X"80",X"E6",X"03",X"C6",X"4C",X"77",X"C9",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"2D",X"24",X"CB",X"FD",X"71",X"24",X"36",X"00",X"24",X"C9",
		X"24",X"2C",X"3A",X"41",X"7A",X"96",X"D6",X"02",X"C6",X"04",X"D0",X"24",X"3A",X"41",X"7B",X"96",
		X"D6",X"02",X"C6",X"04",X"D0",X"2D",X"26",X"7D",X"36",X"30",X"C9",X"24",X"2C",X"3A",X"45",X"7A",
		X"96",X"D6",X"02",X"C6",X"04",X"D0",X"24",X"3A",X"45",X"7B",X"96",X"D6",X"02",X"C6",X"04",X"D0",
		X"2D",X"26",X"7D",X"36",X"30",X"C9",X"16",X"79",X"DD",X"5D",X"EB",X"36",X"02",X"16",X"79",X"DD",
		X"5D",X"EB",X"2C",X"36",X"00",X"2D",X"26",X"7C",X"36",X"3C",X"CB",X"FD",X"36",X"2A",X"24",X"36",
		X"01",X"CB",X"BD",X"24",X"3A",X"A6",X"81",X"77",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",
		X"7F",X"36",X"00",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",X"86",X"31",X"26",
		X"7D",X"CB",X"FD",X"35",X"20",X"3E",X"26",X"79",X"5E",X"2C",X"56",X"2D",X"1A",X"26",X"7D",X"77",
		X"13",X"1A",X"13",X"26",X"79",X"73",X"2C",X"72",X"2D",X"26",X"7B",X"EB",X"21",X"B1",X"2F",X"CD",
		X"83",X"33",X"EB",X"26",X"7D",X"CB",X"BD",X"2C",X"35",X"28",X"03",X"2D",X"18",X"18",X"11",X"47",
		X"2F",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"EB",X"7E",X"FE",X"03",X"CA",
		X"86",X"31",X"18",X"02",X"CB",X"BD",X"26",X"7F",X"7E",X"A7",X"20",X"1A",X"26",X"7A",X"2C",X"3A",
		X"B1",X"81",X"BE",X"38",X"34",X"3A",X"01",X"80",X"E6",X"07",X"20",X"2D",X"2D",X"26",X"7D",X"35",
		X"20",X"27",X"26",X"7F",X"36",X"18",X"35",X"7E",X"FE",X"0C",X"20",X"10",X"E5",X"CD",X"87",X"32",
		X"E1",X"25",X"CD",X"4B",X"0F",X"A6",X"3C",X"25",X"77",X"26",X"7F",X"7E",X"0F",X"0F",X"E6",X"07",
		X"EB",X"21",X"AB",X"2F",X"D7",X"7E",X"16",X"7C",X"12",X"16",X"7C",X"DD",X"5D",X"1C",X"3A",X"1C",
		X"80",X"12",X"16",X"7A",X"1D",X"CD",X"91",X"30",X"C3",X"79",X"30",X"3C",X"3D",X"3E",X"3F",X"3E",
		X"3D",X"00",X"10",X"02",X"10",X"04",X"10",X"06",X"10",X"08",X"10",X"08",X"0E",X"08",X"0C",X"08",
		X"0A",X"08",X"08",X"08",X"06",X"08",X"04",X"08",X"02",X"08",X"00",X"06",X"00",X"04",X"00",X"02",
		X"00",X"00",X"00",X"FE",X"00",X"FC",X"00",X"FA",X"00",X"F8",X"00",X"F8",X"02",X"F8",X"04",X"F8",
		X"06",X"F8",X"08",X"F8",X"0A",X"F8",X"0C",X"F8",X"0E",X"F8",X"10",X"FA",X"10",X"FC",X"10",X"FE",
		X"10",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"66",
		X"21",X"00",X"79",X"11",X"01",X"79",X"01",X"FF",X"06",X"36",X"00",X"ED",X"B0",X"21",X"79",X"30",
		X"22",X"00",X"78",X"22",X"4E",X"78",X"21",X"00",X"78",X"11",X"02",X"78",X"01",X"3E",X"00",X"ED",
		X"B0",X"21",X"4E",X"78",X"11",X"50",X"78",X"01",X"32",X"00",X"ED",X"B0",X"21",X"4E",X"7C",X"11",
		X"50",X"7C",X"01",X"24",X"00",X"36",X"1E",X"ED",X"B0",X"21",X"4F",X"79",X"11",X"50",X"79",X"01",
		X"24",X"00",X"36",X"80",X"2D",X"36",X"00",X"ED",X"B0",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"F7",
		X"3A",X"2A",X"80",X"A7",X"20",X"AA",X"DD",X"E5",X"DD",X"21",X"00",X"78",X"06",X"20",X"CD",X"54",
		X"04",X"DD",X"2C",X"DD",X"2C",X"10",X"F7",X"DD",X"21",X"4E",X"78",X"06",X"19",X"CD",X"54",X"04",
		X"DD",X"2C",X"DD",X"2C",X"10",X"F7",X"DD",X"E1",X"C9",X"F7",X"16",X"7F",X"DD",X"5D",X"EB",X"7E",
		X"A7",X"C8",X"3D",X"21",X"83",X"3C",X"CF",X"7E",X"DD",X"77",X"00",X"23",X"7E",X"DD",X"77",X"01",
		X"C9",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"7C",
		X"1C",X"12",X"14",X"1A",X"67",X"1D",X"1A",X"6F",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",
		X"1C",X"7C",X"12",X"15",X"1A",X"14",X"C6",X"01",X"FE",X"29",X"30",X"06",X"1A",X"FE",X"1F",X"DA",
		X"1D",X"00",X"1D",X"15",X"15",X"EB",X"AF",X"77",X"CB",X"FD",X"77",X"CB",X"BD",X"3E",X"06",X"84",
		X"67",X"36",X"00",X"C9",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"CB",X"FB",X"1A",X"CF",X"CB",X"BB",
		X"7D",X"12",X"1C",X"7C",X"12",X"C3",X"B4",X"30",X"1A",X"6F",X"1C",X"1A",X"67",X"1D",X"3A",X"14",
		X"80",X"ED",X"44",X"CF",X"7D",X"12",X"1C",X"7C",X"12",X"C3",X"B4",X"30",X"1A",X"6F",X"1C",X"1A",
		X"67",X"1D",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"7C",X"1C",X"12",X"14",X"1A",X"67",
		X"1D",X"1A",X"6F",X"CB",X"FB",X"1A",X"CB",X"BB",X"CF",X"7D",X"12",X"1C",X"7C",X"12",X"C9",X"24",
		X"24",X"24",X"2C",X"36",X"07",X"2D",X"24",X"36",X"FF",X"11",X"32",X"31",X"DD",X"73",X"00",X"DD",
		X"72",X"01",X"3E",X"05",X"DD",X"84",X"57",X"DD",X"5D",X"EB",X"34",X"7E",X"FE",X"08",X"20",X"0A",
		X"25",X"25",X"25",X"2C",X"35",X"24",X"34",X"2D",X"24",X"24",X"4F",X"CB",X"3F",X"CB",X"3F",X"FE",
		X"05",X"28",X"26",X"EB",X"21",X"6F",X"31",X"CF",X"15",X"7E",X"12",X"15",X"15",X"15",X"1C",X"23",
		X"79",X"E6",X"03",X"07",X"07",X"86",X"12",X"1D",X"14",X"CD",X"91",X"30",X"C3",X"79",X"30",X"70",
		X"00",X"71",X"00",X"74",X"03",X"78",X"03",X"7C",X"03",X"24",X"24",X"36",X"00",X"3E",X"FA",X"84",
		X"67",X"36",X"00",X"C3",X"79",X"30",X"26",X"7C",X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"11",
		X"98",X"31",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"E6",X"07",X"20",X"2A",X"79",X"0F",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"29",X"FE",X"02",
		X"CC",X"02",X"32",X"FE",X"05",X"CC",X"0C",X"32",X"EB",X"21",X"F4",X"31",X"CF",X"15",X"7E",X"12",
		X"23",X"16",X"79",X"1C",X"7E",X"12",X"1D",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7A",
		X"EB",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"25",X"36",X"A6",X"2C",X"36",X"0D",X"F7",X"16",X"7C",
		X"DD",X"5D",X"3A",X"01",X"80",X"0F",X"0F",X"E6",X"01",X"C6",X"A6",X"12",X"16",X"7A",X"CD",X"E8",
		X"30",X"C3",X"79",X"30",X"60",X"00",X"61",X"00",X"64",X"03",X"68",X"03",X"6C",X"03",X"62",X"00",
		X"63",X"00",X"4C",X"26",X"7A",X"2C",X"35",X"24",X"34",X"2D",X"61",X"C9",X"4C",X"26",X"7A",X"2C",
		X"34",X"24",X"35",X"2D",X"61",X"C9",X"26",X"7C",X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"11",
		X"28",X"32",X"DD",X"73",X"00",X"DD",X"72",X"01",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"E6",X"03",X"20",X"29",X"79",X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"29",X"FE",X"02",X"CC",
		X"02",X"32",X"FE",X"05",X"CC",X"0C",X"32",X"EB",X"21",X"F4",X"31",X"CF",X"15",X"7E",X"12",X"23",
		X"16",X"79",X"1C",X"7E",X"12",X"1D",X"14",X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7A",X"EB",
		X"CD",X"E8",X"30",X"C3",X"79",X"30",X"26",X"7F",X"36",X"00",X"26",X"79",X"36",X"00",X"C3",X"79",
		X"30",X"3A",X"01",X"80",X"E6",X"07",X"C0",X"35",X"C0",X"E5",X"CD",X"87",X"32",X"E1",X"24",X"CD",
		X"4B",X"0F",X"A6",X"25",X"3C",X"77",X"C9",X"48",X"21",X"4E",X"79",X"06",X"13",X"7E",X"3D",X"28",
		X"2A",X"2C",X"2C",X"10",X"F8",X"41",X"C9",X"21",X"4E",X"79",X"06",X"13",X"7E",X"3D",X"28",X"24",
		X"2C",X"2C",X"10",X"F8",X"C9",X"36",X"02",X"16",X"7A",X"DD",X"5D",X"24",X"1A",X"77",X"1C",X"2C",
		X"1A",X"77",X"14",X"24",X"1A",X"77",X"1D",X"2D",X"1A",X"77",X"C9",X"CD",X"A5",X"32",X"CB",X"D4",
		X"36",X"06",X"41",X"C9",X"CD",X"A5",X"32",X"EB",X"CB",X"FB",X"21",X"B3",X"3D",X"79",X"CD",X"83",
		X"33",X"EB",X"CB",X"BD",X"26",X"7F",X"36",X"07",X"C9",X"16",X"7A",X"DD",X"5D",X"1C",X"1A",X"4F",
		X"3A",X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",
		X"D6",X"20",X"0F",X"0F",X"0F",X"E6",X"1F",X"4F",X"C5",X"06",X"05",X"C5",X"CD",X"97",X"32",X"C1",
		X"79",X"C6",X"02",X"E6",X"1F",X"4F",X"10",X"F3",X"C1",X"C9",X"C5",X"01",X"00",X"10",X"C5",X"CD",
		X"97",X"32",X"C1",X"79",X"3C",X"3C",X"E6",X"1E",X"4F",X"10",X"F3",X"21",X"76",X"7A",X"11",X"78",
		X"7A",X"01",X"08",X"00",X"ED",X"B0",X"21",X"76",X"7B",X"11",X"78",X"7B",X"01",X"08",X"00",X"ED",
		X"B0",X"21",X"5D",X"33",X"11",X"F8",X"7A",X"06",X"04",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",
		X"21",X"61",X"33",X"11",X"F8",X"7B",X"06",X"04",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",X"3E",
		X"09",X"06",X"04",X"21",X"78",X"7F",X"77",X"2C",X"2C",X"10",X"FB",X"C1",X"C9",X"20",X"00",X"E0",
		X"00",X"00",X"E0",X"00",X"20",X"E5",X"1A",X"4F",X"3A",X"47",X"7A",X"91",X"6F",X"14",X"1A",X"4F",
		X"3A",X"47",X"7B",X"91",X"67",X"CD",X"B2",X"0E",X"C6",X"04",X"E1",X"CB",X"FB",X"1D",X"0F",X"0F",
		X"0F",X"E6",X"1F",X"CF",X"7E",X"12",X"23",X"15",X"7E",X"12",X"C9",X"CD",X"4B",X"0F",X"E6",X"1F",
		X"FE",X"19",X"30",X"F7",X"C6",X"03",X"77",X"C9",X"E5",X"21",X"47",X"7B",X"CD",X"4B",X"0F",X"E6",
		X"1F",X"FE",X"19",X"30",X"F7",X"C6",X"03",X"5F",X"96",X"D6",X"08",X"C6",X"10",X"7B",X"38",X"EC",
		X"E1",X"77",X"C9",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"2B",X"80",X"A7",X"C8",X"47",X"3A",X"2C",
		X"80",X"21",X"03",X"3C",X"D7",X"11",X"74",X"7F",X"7E",X"12",X"23",X"1C",X"1C",X"10",X"F9",X"C9",
		X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"2D",X"80",X"A7",X"C8",X"21",X"20",X"7F",X"47",X"36",X"01",
		X"2C",X"2C",X"10",X"FA",X"C9",X"F7",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"22",X"84",X"A7",X"C8",
		X"3E",X"3C",X"32",X"23",X"84",X"F7",X"3A",X"2A",X"80",X"A7",X"20",X"E9",X"21",X"23",X"84",X"35",
		X"C0",X"21",X"2D",X"80",X"34",X"21",X"22",X"84",X"35",X"28",X"DA",X"18",X"E3",X"16",X"79",X"DD",
		X"5D",X"EB",X"36",X"02",X"2C",X"36",X"80",X"26",X"7B",X"CD",X"8B",X"33",X"25",X"EB",X"21",X"73",
		X"3D",X"CD",X"65",X"33",X"EB",X"26",X"7C",X"36",X"00",X"F7",X"16",X"79",X"DD",X"5D",X"EB",X"7E",
		X"FE",X"03",X"28",X"1D",X"3A",X"01",X"80",X"0F",X"4F",X"E6",X"03",X"26",X"7C",X"77",X"79",X"0F",
		X"0F",X"E6",X"03",X"C6",X"26",X"2C",X"77",X"2D",X"26",X"7A",X"EB",X"CD",X"91",X"30",X"C3",X"79",
		X"30",X"26",X"7D",X"36",X"FF",X"11",X"5D",X"34",X"26",X"78",X"73",X"2C",X"72",X"16",X"7D",X"DD",
		X"5D",X"EB",X"34",X"7E",X"0F",X"FE",X"04",X"28",X"0D",X"C6",X"04",X"25",X"77",X"26",X"7A",X"EB",
		X"CD",X"91",X"30",X"C3",X"79",X"30",X"26",X"79",X"36",X"00",X"26",X"7F",X"36",X"00",X"C3",X"79",
		X"30",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"34",X"2A",X"1E",X"7A",X"3E",X"10",X"BC",X"28",X"0E",
		X"3E",X"01",X"32",X"07",X"A0",X"3E",X"10",X"CF",X"22",X"1E",X"7A",X"C3",X"47",X"38",X"11",X"A7",
		X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"2F",X"80",X"A7",X"20",X"48",X"3A",X"1C",X"79",
		X"FE",X"03",X"28",X"08",X"3E",X"01",X"32",X"07",X"A0",X"C3",X"47",X"38",X"3E",X"1D",X"32",X"40",
		X"80",X"3E",X"03",X"32",X"1E",X"7D",X"11",X"CF",X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"21",
		X"1E",X"7D",X"35",X"20",X"0E",X"3E",X"06",X"32",X"40",X"80",X"11",X"E3",X"34",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"30",X"BC",X"28",X"30",X"3A",X"14",X"80",X"ED",X"44",
		X"CF",X"22",X"1E",X"7A",X"C9",X"11",X"F5",X"34",X"DD",X"73",X"00",X"DD",X"72",X"01",X"3A",X"1C",
		X"79",X"FE",X"03",X"28",X"B7",X"2A",X"1E",X"7A",X"3E",X"F8",X"BC",X"28",X"0E",X"3E",X"F8",X"CF",
		X"22",X"1E",X"7A",X"3E",X"01",X"32",X"07",X"A0",X"C3",X"47",X"38",X"AF",X"32",X"1E",X"79",X"32",
		X"1E",X"7F",X"C3",X"79",X"30",X"3E",X"02",X"32",X"1C",X"79",X"3E",X"10",X"32",X"1C",X"7C",X"3E",
		X"3C",X"32",X"9C",X"7C",X"2A",X"1E",X"7B",X"22",X"1C",X"7B",X"F7",X"3A",X"1C",X"79",X"FE",X"03",
		X"28",X"29",X"3A",X"1E",X"79",X"3D",X"28",X"1A",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"E6",X"0C",
		X"C6",X"80",X"32",X"1D",X"79",X"2A",X"1E",X"7A",X"22",X"1C",X"7A",X"3A",X"40",X"80",X"32",X"1D",
		X"7C",X"C9",X"32",X"1C",X"79",X"32",X"1C",X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",
		X"37",X"11",X"7A",X"35",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"22",X"1C",X"7A",
		X"2A",X"1E",X"7B",X"22",X"1C",X"7B",X"CD",X"F8",X"37",X"3A",X"1C",X"79",X"FE",X"04",X"C0",X"11",
		X"A5",X"35",X"DD",X"73",X"00",X"DD",X"72",X"01",X"21",X"9C",X"7A",X"36",X"D0",X"24",X"36",X"00",
		X"3E",X"08",X"32",X"1D",X"79",X"3A",X"01",X"80",X"0F",X"4F",X"E6",X"03",X"C6",X"B8",X"32",X"1C",
		X"7C",X"79",X"E6",X"07",X"C6",X"15",X"32",X"1D",X"7C",X"11",X"1C",X"7A",X"CD",X"D4",X"30",X"C3",
		X"79",X"30",X"3E",X"02",X"32",X"1A",X"79",X"AF",X"32",X"1B",X"79",X"3C",X"32",X"1A",X"7D",X"3E",
		X"5C",X"32",X"1A",X"7C",X"3E",X"30",X"32",X"9A",X"7C",X"2A",X"1E",X"7B",X"3E",X"02",X"84",X"67",
		X"22",X"1A",X"7B",X"3A",X"A7",X"81",X"32",X"1A",X"7E",X"F7",X"3A",X"1A",X"79",X"FE",X"03",X"28",
		X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",X"1E",
		X"7A",X"3E",X"FE",X"84",X"67",X"22",X"1A",X"7A",X"3A",X"40",X"80",X"32",X"1B",X"7C",X"21",X"1A",
		X"7D",X"CD",X"71",X"32",X"C9",X"32",X"1A",X"79",X"32",X"1A",X"7F",X"C3",X"79",X"30",X"DD",X"5D",
		X"6B",X"CD",X"EE",X"37",X"11",X"2D",X"36",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",
		X"3E",X"FE",X"84",X"67",X"22",X"1A",X"7A",X"2A",X"1E",X"7B",X"3E",X"02",X"84",X"67",X"22",X"1A",
		X"7B",X"CD",X"F8",X"37",X"3A",X"1A",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"3E",X"02",X"32",
		X"18",X"79",X"AF",X"32",X"19",X"79",X"3C",X"32",X"18",X"7D",X"3E",X"5D",X"32",X"18",X"7C",X"3E",
		X"30",X"32",X"98",X"7C",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",X"18",X"7B",X"3A",X"A7",
		X"81",X"32",X"18",X"7E",X"F7",X"3A",X"18",X"79",X"FE",X"03",X"28",X"2D",X"3A",X"1C",X"79",X"FE",
		X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",X"1E",X"7A",X"3E",X"FE",X"84",X"67",
		X"22",X"18",X"7A",X"3A",X"40",X"80",X"32",X"19",X"7C",X"21",X"18",X"7D",X"CD",X"71",X"32",X"C9",
		X"32",X"18",X"79",X"32",X"18",X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",X"37",X"11",
		X"B8",X"36",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"FE",X"84",X"67",X"22",
		X"18",X"7A",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",X"18",X"7B",X"CD",X"F8",X"37",X"3A",
		X"18",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"3E",X"02",X"32",X"16",X"79",X"AF",X"32",X"17",
		X"79",X"3C",X"32",X"16",X"7D",X"3E",X"5E",X"32",X"16",X"7C",X"3E",X"30",X"32",X"96",X"7C",X"2A",
		X"1E",X"7B",X"3E",X"02",X"84",X"67",X"22",X"16",X"7B",X"3A",X"A7",X"81",X"32",X"16",X"7E",X"F7",
		X"3A",X"16",X"79",X"FE",X"03",X"28",X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",
		X"79",X"3D",X"28",X"17",X"2A",X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"16",X"7A",X"3A",X"40",
		X"80",X"32",X"17",X"7C",X"21",X"16",X"7D",X"CD",X"71",X"32",X"C9",X"32",X"16",X"79",X"32",X"16",
		X"7F",X"C3",X"79",X"30",X"DD",X"5D",X"6B",X"CD",X"EE",X"37",X"11",X"43",X"37",X"DD",X"73",X"00",
		X"DD",X"72",X"01",X"2A",X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"16",X"7A",X"2A",X"1E",X"7B",
		X"3E",X"02",X"84",X"67",X"22",X"16",X"7B",X"CD",X"F8",X"37",X"3A",X"16",X"79",X"FE",X"04",X"C0",
		X"AF",X"18",X"C8",X"3E",X"02",X"32",X"14",X"79",X"AF",X"32",X"15",X"79",X"3C",X"32",X"14",X"7D",
		X"3E",X"5F",X"32",X"14",X"7C",X"3E",X"30",X"32",X"94",X"7C",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",
		X"67",X"22",X"14",X"7B",X"3A",X"A7",X"81",X"32",X"14",X"7E",X"F7",X"3A",X"14",X"79",X"FE",X"03",
		X"28",X"2D",X"3A",X"1C",X"79",X"FE",X"03",X"28",X"26",X"3A",X"1E",X"79",X"3D",X"28",X"17",X"2A",
		X"1E",X"7A",X"3E",X"02",X"84",X"67",X"22",X"14",X"7A",X"3A",X"40",X"80",X"32",X"15",X"7C",X"21",
		X"14",X"7D",X"CD",X"71",X"32",X"C9",X"32",X"14",X"79",X"32",X"14",X"7F",X"C3",X"79",X"30",X"DD",
		X"5D",X"6B",X"CD",X"EE",X"37",X"11",X"CE",X"37",X"DD",X"73",X"00",X"DD",X"72",X"01",X"2A",X"1E",
		X"7A",X"3E",X"02",X"84",X"67",X"22",X"14",X"7A",X"2A",X"1E",X"7B",X"3E",X"FE",X"84",X"67",X"22",
		X"14",X"7B",X"CD",X"F8",X"37",X"3A",X"14",X"79",X"FE",X"04",X"C0",X"AF",X"18",X"C8",X"26",X"7C",
		X"2C",X"36",X"0C",X"2D",X"24",X"36",X"FF",X"C9",X"16",X"7D",X"DD",X"5D",X"EB",X"34",X"7E",X"4F",
		X"0F",X"0F",X"E6",X"07",X"D6",X"05",X"C6",X"03",X"DC",X"3D",X"38",X"79",X"E6",X"03",X"C0",X"79",
		X"0F",X"0F",X"E6",X"07",X"FE",X"07",X"28",X"0F",X"EB",X"21",X"2F",X"38",X"CF",X"15",X"7E",X"12",
		X"23",X"1C",X"16",X"79",X"7E",X"12",X"C9",X"25",X"36",X"00",X"26",X"79",X"36",X"04",X"C9",X"60",
		X"00",X"61",X"00",X"64",X"03",X"68",X"03",X"6C",X"03",X"62",X"00",X"63",X"00",X"26",X"7A",X"2C",
		X"35",X"24",X"34",X"2D",X"26",X"7D",X"C9",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"E6",X"07",X"21",
		X"58",X"38",X"D7",X"7E",X"32",X"40",X"80",X"C9",X"02",X"03",X"04",X"05",X"06",X"05",X"04",X"03",
		X"3E",X"03",X"32",X"12",X"79",X"32",X"13",X"79",X"3E",X"58",X"32",X"12",X"7C",X"2A",X"1E",X"7B",
		X"3E",X"05",X"84",X"67",X"22",X"12",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"FB",X"84",X"67",X"22",
		X"12",X"7A",X"3A",X"40",X"80",X"32",X"13",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",
		X"12",X"79",X"32",X"12",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"10",X"79",X"32",X"11",X"79",
		X"3E",X"80",X"32",X"10",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"10",X"7B",X"F7",X"2A",X"1E",X"7A",
		X"3E",X"FB",X"84",X"67",X"22",X"10",X"7A",X"3A",X"40",X"80",X"32",X"11",X"7C",X"3A",X"1E",X"79",
		X"FE",X"01",X"C0",X"AF",X"32",X"10",X"79",X"32",X"10",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",
		X"0E",X"79",X"32",X"0F",X"79",X"3E",X"84",X"32",X"0E",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",X"84",
		X"67",X"22",X"0E",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"FB",X"84",X"67",X"22",X"0E",X"7A",X"3A",
		X"40",X"80",X"32",X"0F",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"0E",X"79",X"32",
		X"0E",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"0C",X"79",X"32",X"0D",X"79",X"3E",X"88",X"32",
		X"0C",X"7C",X"2A",X"1E",X"7B",X"3E",X"05",X"84",X"67",X"22",X"0C",X"7B",X"F7",X"2A",X"1E",X"7A",
		X"25",X"22",X"0C",X"7A",X"3A",X"40",X"80",X"32",X"0D",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",
		X"AF",X"32",X"0C",X"79",X"32",X"0C",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"0A",X"79",X"32",
		X"0B",X"79",X"3E",X"8C",X"32",X"0A",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"0A",X"7B",X"F7",X"2A",
		X"1E",X"7A",X"25",X"22",X"0A",X"7A",X"3A",X"40",X"80",X"32",X"0B",X"7C",X"3A",X"1E",X"79",X"FE",
		X"01",X"C0",X"AF",X"32",X"0A",X"79",X"32",X"0A",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"08",
		X"79",X"32",X"09",X"79",X"3E",X"90",X"32",X"08",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",X"84",X"67",
		X"22",X"08",X"7B",X"F7",X"2A",X"1E",X"7A",X"25",X"22",X"08",X"7A",X"3A",X"40",X"80",X"32",X"09",
		X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"08",X"79",X"32",X"08",X"7F",X"C3",X"79",
		X"30",X"3E",X"03",X"32",X"06",X"79",X"32",X"07",X"79",X"3E",X"94",X"32",X"06",X"7C",X"2A",X"1E",
		X"7B",X"3E",X"05",X"84",X"67",X"22",X"06",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"03",X"84",X"67",
		X"22",X"06",X"7A",X"3A",X"40",X"80",X"32",X"07",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",
		X"32",X"06",X"79",X"32",X"06",X"7F",X"C3",X"79",X"30",X"3E",X"03",X"32",X"04",X"79",X"32",X"05",
		X"79",X"3E",X"98",X"32",X"04",X"7C",X"2A",X"1E",X"7B",X"24",X"22",X"04",X"7B",X"F7",X"2A",X"1E",
		X"7A",X"3E",X"03",X"84",X"67",X"22",X"04",X"7A",X"3A",X"40",X"80",X"32",X"05",X"7C",X"3A",X"1E",
		X"79",X"FE",X"01",X"C0",X"AF",X"32",X"04",X"79",X"32",X"04",X"7F",X"C3",X"79",X"30",X"3E",X"03",
		X"32",X"02",X"79",X"32",X"03",X"79",X"3E",X"9C",X"32",X"02",X"7C",X"2A",X"1E",X"7B",X"3E",X"FD",
		X"84",X"67",X"22",X"02",X"7B",X"F7",X"2A",X"1E",X"7A",X"3E",X"03",X"84",X"67",X"22",X"02",X"7A",
		X"3A",X"40",X"80",X"32",X"03",X"7C",X"3A",X"1E",X"79",X"FE",X"01",X"C0",X"AF",X"32",X"02",X"79",
		X"32",X"02",X"7F",X"C3",X"79",X"30",X"3A",X"28",X"80",X"A7",X"20",X"59",X"16",X"79",X"DD",X"5D",
		X"EB",X"36",X"02",X"2C",X"36",X"00",X"26",X"7C",X"2D",X"36",X"00",X"11",X"64",X"3A",X"DD",X"73",
		X"00",X"DD",X"72",X"01",X"16",X"79",X"DD",X"5D",X"1A",X"FE",X"03",X"28",X"08",X"16",X"7A",X"CD",
		X"E8",X"30",X"C3",X"79",X"30",X"16",X"7D",X"3E",X"80",X"12",X"21",X"CD",X"3E",X"11",X"B6",X"3A",
		X"C5",X"06",X"13",X"1A",X"0F",X"BE",X"20",X"29",X"13",X"23",X"10",X"F7",X"CD",X"C9",X"3A",X"11",
		X"99",X"3A",X"DD",X"73",X"00",X"DD",X"72",X"01",X"C1",X"16",X"7D",X"DD",X"5D",X"EB",X"35",X"C0",
		X"C5",X"CD",X"7C",X"3B",X"C1",X"16",X"79",X"DD",X"5D",X"AF",X"12",X"16",X"7F",X"12",X"C3",X"79",
		X"30",X"CD",X"09",X"3B",X"18",X"D9",X"5A",X"5C",X"50",X"48",X"02",X"12",X"10",X"04",X"48",X"2E",
		X"14",X"2C",X"18",X"30",X"48",X"2A",X"3A",X"1A",X"A0",X"21",X"E1",X"3A",X"CD",X"48",X"3B",X"21",
		X"21",X"19",X"06",X"07",X"0E",X"B0",X"3E",X"1A",X"CD",X"5D",X"14",X"21",X"F1",X"3A",X"C3",X"62",
		X"3B",X"D0",X"CF",X"CE",X"CD",X"CC",X"CB",X"CA",X"DB",X"E7",X"E4",X"ED",X"EF",X"ED",X"E8",X"F5",
		X"EA",X"DB",X"DB",X"DB",X"DB",X"DB",X"BA",X"B8",X"BB",X"C3",X"B8",X"C9",X"BD",X"DB",X"C8",X"B1",
		X"DB",X"F1",X"E0",X"F1",X"DC",X"E7",X"E7",X"DB",X"DB",X"21",X"20",X"3B",X"CD",X"48",X"3B",X"21",
		X"21",X"19",X"06",X"09",X"0E",X"B0",X"3E",X"1B",X"CD",X"5D",X"14",X"21",X"30",X"3B",X"18",X"42",
		X"F2",X"F1",X"F5",X"F2",X"DB",X"F3",X"E7",X"E6",X"DD",X"DB",X"E9",X"F5",X"EB",X"ED",X"E8",X"EF",
		X"C7",X"BB",X"BA",X"B1",X"DB",X"B5",X"BC",X"C6",X"C5",X"B8",X"DB",X"E8",X"F5",X"E9",X"F3",X"E7",
		X"DB",X"BA",X"B8",X"BB",X"C3",X"B8",X"C9",X"BD",X"11",X"80",X"84",X"06",X"10",X"7E",X"2F",X"12",
		X"23",X"13",X"10",X"F9",X"21",X"21",X"19",X"11",X"80",X"84",X"06",X"10",X"0E",X"C0",X"CD",X"1F",
		X"14",X"C9",X"11",X"80",X"84",X"06",X"18",X"7E",X"2F",X"12",X"23",X"13",X"10",X"F9",X"21",X"22",
		X"17",X"11",X"80",X"84",X"06",X"18",X"0E",X"C0",X"CD",X"1F",X"14",X"C9",X"21",X"21",X"19",X"06",
		X"10",X"0E",X"C0",X"3E",X"24",X"CD",X"5D",X"14",X"21",X"21",X"19",X"06",X"10",X"0E",X"B0",X"3E",
		X"24",X"CD",X"5D",X"14",X"21",X"22",X"17",X"06",X"18",X"0E",X"C0",X"C3",X"5D",X"14",X"21",X"00",
		X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",X"21",X"01",X"3C",X"01",X"01",X"64",X"CD",X"10",
		X"01",X"F7",X"21",X"60",X"80",X"01",X"04",X"74",X"CD",X"E5",X"00",X"F7",X"3A",X"63",X"80",X"FE",
		X"05",X"C2",X"00",X"00",X"F7",X"21",X"02",X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",X"21",
		X"60",X"80",X"01",X"04",X"74",X"CD",X"E5",X"00",X"F7",X"3A",X"63",X"80",X"FE",X"95",X"C2",X"00",
		X"00",X"F7",X"C9",X"21",X"9E",X"3B",X"11",X"F6",X"3B",X"06",X"0A",X"1A",X"BE",X"C2",X"00",X"00",
		X"23",X"13",X"10",X"F7",X"F7",X"C9",X"21",X"00",X"3C",X"01",X"01",X"64",X"CD",X"10",X"01",X"F7",
		X"10",X"80",X"E5",X"00",X"0A",X"0A",X"0A",X"0A",X"0A",X"0A",X"0B",X"0B",X"0B",X"0B",X"0B",X"0B",
		X"55",X"55",X"55",X"55",X"55",X"55",X"56",X"56",X"56",X"56",X"56",X"56",X"0F",X"0F",X"0F",X"0F",
		X"0F",X"0F",X"0C",X"0C",X"0C",X"0C",X"0C",X"0C",X"0B",X"0B",X"08",X"08",X"08",X"08",X"08",X"08",
		X"0D",X"0D",X"0D",X"0D",X"0D",X"0D",X"0E",X"0E",X"0E",X"12",X"12",X"12",X"13",X"13",X"13",X"14",
		X"14",X"14",X"14",X"14",X"14",X"0E",X"0E",X"0E",X"10",X"10",X"10",X"10",X"10",X"10",X"14",X"14",
		X"14",X"11",X"11",X"11",X"11",X"11",X"11",X"16",X"16",X"16",X"16",X"17",X"17",X"17",X"17",X"0F",
		X"0F",X"08",X"08",X"08",X"08",X"55",X"55",X"10",X"10",X"08",X"08",X"08",X"08",X"11",X"11",X"14",
		X"14",X"15",X"15",X"15",X"15",X"08",X"08",X"08",X"08",X"0E",X"0E",X"78",X"79",X"7A",X"7B",X"7C",
		X"7D",X"7E",X"7F",X"23",X"2B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"6D",X"2B",X"79",
		X"2B",X"0D",X"34",X"F8",X"1E",X"00",X"20",X"18",X"20",X"36",X"22",X"C4",X"21",X"B1",X"21",X"E7",
		X"20",X"A8",X"23",X"87",X"24",X"67",X"25",X"D7",X"25",X"2E",X"26",X"84",X"26",X"DF",X"26",X"36",
		X"27",X"4C",X"28",X"45",X"1B",X"18",X"1C",X"00",X"1C",X"0C",X"1C",X"61",X"1E",X"60",X"1A",X"F0",
		X"1A",X"89",X"1A",X"61",X"1C",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2D",X"1B",X"39",
		X"1B",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"83",X"2B",X"DE",X"1C",X"D6",X"2E",X"00",
		X"00",X"00",X"00",X"DD",X"28",X"2E",X"2A",X"00",X"00",X"00",X"00",X"96",X"2B",X"A6",X"2B",X"E4",
		X"2B",X"2E",X"2C",X"77",X"2C",X"C4",X"2C",X"10",X"2D",X"5C",X"2D",X"A3",X"2D",X"B7",X"2D",X"C8",
		X"2D",X"F9",X"2D",X"60",X"38",X"98",X"38",X"CD",X"38",X"05",X"39",X"3A",X"39",X"6C",X"39",X"A1",
		X"39",X"D9",X"39",X"0E",X"3A",X"25",X"35",X"81",X"34",X"00",X"00",X"00",X"00",X"00",X"00",X"C2",
		X"35",X"4D",X"36",X"D8",X"36",X"63",X"37",X"46",X"3A",X"5C",X"1F",X"06",X"23",X"AC",X"22",X"00",
		X"00",X"01",X"00",X"00",X"02",X"00",X"00",X"03",X"00",X"00",X"05",X"00",X"00",X"07",X"00",X"00",
		X"10",X"00",X"00",X"15",X"00",X"00",X"20",X"00",X"00",X"25",X"00",X"00",X"30",X"00",X"00",X"40",
		X"00",X"00",X"50",X"00",X"00",X"60",X"00",X"00",X"70",X"00",X"00",X"80",X"00",X"00",X"90",X"00",
		X"00",X"00",X"01",X"00",X"50",X"01",X"00",X"00",X"02",X"00",X"50",X"02",X"00",X"00",X"04",X"00",
		X"00",X"10",X"00",X"00",X"40",X"0C",X"3F",X"18",X"3B",X"24",X"35",X"2D",X"2D",X"35",X"24",X"3B",
		X"18",X"3F",X"0C",X"40",X"00",X"3F",X"F4",X"3B",X"E8",X"35",X"DC",X"2D",X"D3",X"24",X"CB",X"18",
		X"C5",X"0C",X"C1",X"00",X"C0",X"F4",X"C1",X"E8",X"C5",X"DC",X"CB",X"D3",X"D3",X"CB",X"DC",X"C5",
		X"E8",X"C1",X"F4",X"C0",X"00",X"C1",X"0C",X"C5",X"18",X"CB",X"24",X"D3",X"2D",X"DC",X"35",X"E8",
		X"3B",X"F4",X"3F",X"00",X"30",X"09",X"2F",X"12",X"2C",X"1B",X"28",X"22",X"22",X"28",X"1B",X"2C",
		X"12",X"2F",X"09",X"30",X"00",X"2F",X"F7",X"2C",X"EE",X"28",X"E5",X"22",X"DE",X"1B",X"D8",X"12",
		X"D4",X"09",X"D1",X"00",X"D0",X"F7",X"D1",X"EE",X"D4",X"E5",X"D8",X"DE",X"DE",X"D8",X"E5",X"D4",
		X"EE",X"D1",X"F7",X"D0",X"00",X"D1",X"09",X"D4",X"12",X"D8",X"1B",X"DE",X"22",X"E5",X"28",X"EE",
		X"2C",X"F7",X"2F",X"00",X"20",X"06",X"1F",X"0C",X"1E",X"11",X"1B",X"17",X"17",X"1B",X"11",X"1E",
		X"0C",X"1F",X"06",X"20",X"00",X"1F",X"FA",X"1E",X"F4",X"1B",X"EF",X"17",X"E9",X"11",X"E5",X"0C",
		X"E2",X"06",X"E1",X"00",X"E0",X"FA",X"E1",X"F4",X"E2",X"EF",X"E5",X"E9",X"E9",X"E5",X"EF",X"E2",
		X"F4",X"E1",X"FA",X"E0",X"00",X"E1",X"06",X"E2",X"0C",X"E5",X"11",X"E9",X"17",X"EF",X"1B",X"F4",
		X"1E",X"FA",X"1F",X"00",X"18",X"05",X"18",X"09",X"16",X"0D",X"14",X"11",X"11",X"14",X"0D",X"16",
		X"09",X"18",X"05",X"18",X"00",X"18",X"FB",X"16",X"F7",X"14",X"F3",X"11",X"EF",X"0D",X"EC",X"09",
		X"EA",X"05",X"E8",X"00",X"E8",X"FB",X"E8",X"F7",X"EA",X"F3",X"EC",X"EF",X"EF",X"EC",X"F3",X"EA",
		X"F7",X"E8",X"FB",X"E8",X"00",X"E8",X"05",X"EA",X"09",X"EC",X"0D",X"EF",X"11",X"F3",X"14",X"F7",
		X"16",X"FB",X"18",X"00",X"10",X"03",X"10",X"06",X"0F",X"09",X"0D",X"0B",X"0B",X"0D",X"09",X"0F",
		X"06",X"10",X"03",X"10",X"00",X"10",X"FD",X"0F",X"FA",X"0D",X"F7",X"0B",X"F5",X"09",X"F3",X"06",
		X"F1",X"03",X"F0",X"00",X"F0",X"FD",X"F0",X"FA",X"F1",X"F7",X"F3",X"F5",X"F5",X"F3",X"F7",X"F1",
		X"FA",X"F0",X"FD",X"F0",X"00",X"F0",X"03",X"F1",X"06",X"F3",X"09",X"F5",X"0B",X"F7",X"0D",X"FA",
		X"0F",X"FD",X"10",X"24",X"00",X"54",X"0E",X"40",X"1A",X"64",X"04",X"2A",X"5C",X"0E",X"04",X"38",
		X"54",X"1A",X"00",X"11",X"12",X"10",X"11",X"24",X"1C",X"0C",X"18",X"1B",X"0E",X"2D",X"2E",X"28",
		X"24",X"01",X"09",X"08",X"02",X"24",X"17",X"0A",X"16",X"0C",X"18",X"24",X"15",X"1D",X"0D",X"50",
		X"2F",X"30",X"31",X"32",X"33",X"34",X"35",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"35");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
