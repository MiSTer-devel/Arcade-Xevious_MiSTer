library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity xevious_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of xevious_cpu2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"C3",X"65",X"01",X"12",X"42",X"21",X"00",X"00",X"87",X"D2",X"58",X"00",X"25",X"C3",X"58",X"00",
		X"A7",X"F2",X"58",X"00",X"25",X"C3",X"58",X"00",X"A7",X"F0",X"ED",X"44",X"C9",X"33",X"33",X"C9",
		X"EB",X"CD",X"05",X"00",X"29",X"19",X"C9",X"FF",X"EB",X"CD",X"05",X"00",X"29",X"29",X"19",X"C9",
		X"E1",X"DD",X"75",X"00",X"DD",X"74",X"01",X"C9",X"3A",X"03",X"80",X"A7",X"3E",X"03",X"28",X"04",
		X"25",X"25",X"3E",X"19",X"85",X"E6",X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",X"67",X"E6",X"C0",
		X"B5",X"6F",X"7C",X"E6",X"07",X"81",X"67",X"C9",X"85",X"6F",X"D0",X"24",X"C9",X"0E",X"12",X"1B",
		X"1B",X"22",X"24",X"16",X"18",X"1E",X"ED",X"45",X"11",X"17",X"93",X"21",X"16",X"93",X"01",X"13",
		X"00",X"ED",X"B8",X"DD",X"21",X"60",X"01",X"1E",X"00",X"01",X"04",X"05",X"DD",X"7E",X"00",X"DD",
		X"23",X"6F",X"26",X"20",X"7E",X"7B",X"81",X"5F",X"7E",X"12",X"10",X"F0",X"06",X"05",X"21",X"04",
		X"93",X"7E",X"2C",X"B6",X"2C",X"2F",X"A6",X"2C",X"A6",X"2C",X"E6",X"0F",X"20",X"04",X"10",X"F1",
		X"18",X"40",X"05",X"28",X"4F",X"05",X"CB",X"20",X"CB",X"20",X"0F",X"38",X"03",X"04",X"18",X"FA",
		X"3A",X"00",X"93",X"CB",X"3F",X"5F",X"CB",X"11",X"C6",X"01",X"6F",X"26",X"93",X"7E",X"CB",X"41",
		X"28",X"04",X"07",X"07",X"07",X"07",X"E6",X"F0",X"B0",X"CB",X"41",X"28",X"04",X"07",X"07",X"07",
		X"07",X"77",X"3A",X"00",X"93",X"A7",X"20",X"02",X"3E",X"02",X"3D",X"32",X"00",X"93",X"7B",X"A7",
		X"28",X"09",X"2A",X"02",X"93",X"7E",X"32",X"01",X"93",X"18",X"42",X"2A",X"02",X"93",X"3A",X"01",
		X"93",X"77",X"18",X"39",X"4F",X"21",X"00",X"93",X"CB",X"41",X"20",X"2D",X"7E",X"CB",X"3F",X"28",
		X"13",X"CB",X"59",X"20",X"0C",X"7E",X"FE",X"05",X"30",X"03",X"34",X"18",X"D5",X"36",X"05",X"18",
		X"D1",X"35",X"18",X"CE",X"2A",X"02",X"93",X"CB",X"59",X"20",X"03",X"2B",X"18",X"01",X"23",X"22",
		X"02",X"93",X"3E",X"01",X"32",X"00",X"93",X"18",X"B9",X"36",X"05",X"18",X"B5",X"21",X"E2",X"C0",
		X"11",X"01",X"93",X"06",X"03",X"1A",X"1C",X"CD",X"51",X"01",X"10",X"F9",X"21",X"E2",X"B0",X"3A",
		X"00",X"93",X"06",X"06",X"A7",X"0E",X"04",X"28",X"02",X"0E",X"0C",X"71",X"2D",X"3D",X"10",X"F4",
		X"C9",X"4F",X"E6",X"0F",X"77",X"2D",X"79",X"07",X"07",X"07",X"07",X"E6",X"0F",X"77",X"2D",X"C9",
		X"FD",X"FB",X"F7",X"EF",X"FE",X"3A",X"09",X"04",X"32",X"72",X"85",X"3A",X"FB",X"15",X"32",X"73",
		X"85",X"31",X"80",X"97",X"21",X"00",X"10",X"11",X"00",X"A4",X"01",X"20",X"00",X"ED",X"B0",X"21",
		X"B6",X"01",X"11",X"C0",X"82",X"01",X"40",X"00",X"ED",X"B0",X"21",X"02",X"80",X"7E",X"3D",X"20",
		X"FC",X"77",X"32",X"0A",X"80",X"3A",X"16",X"80",X"CB",X"7F",X"28",X"EE",X"DD",X"21",X"C0",X"82",
		X"06",X"20",X"C5",X"CD",X"AF",X"01",X"C1",X"DD",X"23",X"DD",X"23",X"10",X"F5",X"18",X"DB",X"DD",
		X"6E",X"00",X"DD",X"66",X"01",X"E9",X"F6",X"01",X"18",X"02",X"8F",X"06",X"8B",X"07",X"27",X"02",
		X"64",X"02",X"CD",X"07",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",X"1F",X"00",
		X"1F",X"00",X"A6",X"02",X"1E",X"03",X"21",X"40",X"82",X"11",X"C0",X"87",X"01",X"40",X"00",X"ED",
		X"B0",X"21",X"40",X"83",X"11",X"C0",X"97",X"01",X"40",X"00",X"ED",X"B0",X"21",X"40",X"81",X"11",
		X"C0",X"A7",X"01",X"40",X"00",X"ED",X"B0",X"C9",X"2A",X"0C",X"80",X"7D",X"6C",X"26",X"D0",X"77",
		X"3A",X"0E",X"80",X"32",X"20",X"D0",X"C9",X"3A",X"18",X"80",X"4F",X"3A",X"29",X"80",X"47",X"91",
		X"C8",X"30",X"1B",X"79",X"32",X"29",X"80",X"FE",X"A0",X"C8",X"90",X"27",X"21",X"00",X"A0",X"86",
		X"27",X"77",X"21",X"5D",X"02",X"11",X"80",X"80",X"01",X"07",X"00",X"ED",X"B0",X"C9",X"27",X"3D",
		X"32",X"22",X"80",X"79",X"32",X"29",X"80",X"3E",X"01",X"32",X"1B",X"80",X"C9",X"30",X"10",X"00",
		X"80",X"FF",X"10",X"10",X"3A",X"2A",X"80",X"A7",X"C0",X"3A",X"01",X"80",X"1F",X"E6",X"03",X"C6",
		X"25",X"21",X"4F",X"7C",X"06",X"13",X"77",X"2C",X"2C",X"10",X"FB",X"3A",X"01",X"80",X"0F",X"0F",
		X"0F",X"E6",X"07",X"4F",X"21",X"96",X"02",X"D7",X"7E",X"32",X"1C",X"80",X"79",X"21",X"9E",X"02",
		X"D7",X"7E",X"32",X"43",X"80",X"C9",X"07",X"08",X"09",X"0A",X"0B",X"0A",X"09",X"08",X"10",X"11",
		X"12",X"13",X"14",X"13",X"12",X"11",X"3A",X"2A",X"80",X"A7",X"C0",X"CD",X"D4",X"02",X"3A",X"03",
		X"80",X"A7",X"3E",X"40",X"28",X"02",X"3E",X"30",X"2A",X"10",X"80",X"CF",X"29",X"29",X"AF",X"29",
		X"17",X"6C",X"67",X"22",X"0C",X"80",X"3A",X"03",X"80",X"A7",X"3E",X"00",X"28",X"02",X"3E",X"00",
		X"32",X"0E",X"80",X"C9",X"2A",X"10",X"80",X"4C",X"3A",X"14",X"80",X"CF",X"22",X"10",X"80",X"3A",
		X"0F",X"80",X"A7",X"C0",X"7C",X"B9",X"C8",X"FA",X"EC",X"02",X"C6",X"40",X"C6",X"F2",X"6F",X"3A",
		X"03",X"80",X"A7",X"3A",X"13",X"80",X"28",X"02",X"C6",X"FE",X"C6",X"FF",X"67",X"01",X"B8",X"20",
		X"16",X"FE",X"5D",X"22",X"00",X"F0",X"EB",X"E5",X"CD",X"38",X"00",X"3A",X"00",X"F0",X"77",X"3E",
		X"10",X"84",X"67",X"3A",X"01",X"F0",X"77",X"E1",X"EB",X"14",X"24",X"10",X"E5",X"C9",X"21",X"00",
		X"79",X"11",X"00",X"83",X"06",X"40",X"E5",X"CD",X"32",X"03",X"E1",X"2C",X"2C",X"1C",X"1C",X"10",
		X"F5",X"C9",X"7E",X"3D",X"C8",X"E5",X"3C",X"20",X"0C",X"4C",X"24",X"77",X"2C",X"77",X"24",X"77",
		X"2D",X"77",X"3C",X"61",X"77",X"2C",X"4E",X"79",X"12",X"D5",X"24",X"56",X"2D",X"5E",X"EB",X"CD",
		X"B3",X"03",X"FE",X"02",X"38",X"03",X"21",X"00",X"00",X"CD",X"89",X"03",X"E5",X"EB",X"24",X"5E",
		X"2C",X"56",X"EB",X"CD",X"B3",X"03",X"A7",X"28",X"02",X"2E",X"00",X"CD",X"A2",X"03",X"D1",X"E1",
		X"2C",X"72",X"25",X"73",X"2D",X"77",X"25",X"EB",X"E1",X"4C",X"24",X"24",X"24",X"7E",X"12",X"2C",
		X"1C",X"7E",X"12",X"61",X"2D",X"14",X"14",X"1D",X"C9",X"3A",X"03",X"80",X"A7",X"28",X"0F",X"3E",
		X"48",X"CB",X"41",X"20",X"02",X"3E",X"58",X"95",X"6F",X"3E",X"01",X"9C",X"67",X"C9",X"3E",X"08",
		X"D7",X"C9",X"3A",X"03",X"80",X"A7",X"3E",X"EF",X"28",X"07",X"85",X"CB",X"49",X"C0",X"C6",X"10",
		X"C9",X"95",X"C9",X"AF",X"29",X"17",X"29",X"17",X"29",X"17",X"6C",X"67",X"C9",X"0A",X"03",X"21",
		X"D8",X"04",X"CF",X"7E",X"32",X"2B",X"80",X"23",X"7E",X"32",X"2C",X"80",X"ED",X"43",X"85",X"81",
		X"C9",X"3A",X"16",X"80",X"2F",X"07",X"07",X"07",X"E6",X"03",X"21",X"08",X"04",X"D7",X"7E",X"6F",
		X"3A",X"88",X"81",X"85",X"FE",X"80",X"38",X"02",X"D6",X"40",X"32",X"88",X"81",X"18",X"D0",X"21",
		X"88",X"81",X"0A",X"86",X"03",X"FE",X"80",X"38",X"02",X"D6",X"40",X"18",X"C2",X"21",X"00",X"00",
		X"22",X"2B",X"80",X"ED",X"43",X"85",X"81",X"C9",X"02",X"00",X"06",X"10",X"ED",X"43",X"85",X"81",
		X"2A",X"81",X"81",X"3A",X"8B",X"81",X"CD",X"2C",X"04",X"11",X"10",X"00",X"A7",X"ED",X"52",X"19",
		X"38",X"02",X"2E",X"10",X"3A",X"88",X"81",X"85",X"32",X"88",X"81",X"C9",X"C5",X"4F",X"AF",X"06",
		X"10",X"29",X"17",X"38",X"03",X"B9",X"38",X"02",X"91",X"23",X"10",X"F5",X"C1",X"C9",X"0A",X"32",
		X"A0",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A3",X"81",X"03",X"ED",X"43",X"85",
		X"81",X"C9",X"0A",X"32",X"A4",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A2",X"81",
		X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A1",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",
		X"0A",X"32",X"A5",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"A6",X"81",X"03",X"ED",
		X"43",X"85",X"81",X"C9",X"0A",X"32",X"A7",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",
		X"B1",X"81",X"03",X"ED",X"43",X"85",X"81",X"C9",X"04",X"0B",X"05",X"0A",X"06",X"09",X"06",X"25",
		X"06",X"5C",X"06",X"29",X"06",X"5E",X"06",X"64",X"06",X"66",X"06",X"72",X"04",X"30",X"04",X"31",
		X"05",X"30",X"06",X"30",X"06",X"3F",X"06",X"48",X"06",X"4B",X"02",X"54",X"03",X"54",X"04",X"54",
		X"02",X"58",X"03",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",
		X"04",X"58",X"04",X"58",X"04",X"58",X"04",X"58",X"03",X"01",X"03",X"01",X"03",X"01",X"04",X"01",
		X"04",X"01",X"04",X"01",X"05",X"01",X"05",X"01",X"05",X"01",X"02",X"19",X"02",X"19",X"02",X"19",
		X"04",X"01",X"04",X"01",X"04",X"04",X"04",X"04",X"04",X"05",X"04",X"05",X"05",X"05",X"05",X"05",
		X"06",X"05",X"06",X"05",X"03",X"19",X"03",X"19",X"04",X"19",X"04",X"19",X"05",X"19",X"05",X"19",
		X"03",X"27",X"03",X"27",X"04",X"27",X"04",X"27",X"05",X"27",X"05",X"27",X"03",X"1F",X"03",X"1F",
		X"04",X"1F",X"04",X"1F",X"05",X"1F",X"05",X"1F",X"03",X"13",X"03",X"13",X"04",X"13",X"04",X"13",
		X"05",X"13",X"05",X"13",X"03",X"36",X"03",X"36",X"03",X"37",X"03",X"37",X"04",X"37",X"04",X"37",
		X"03",X"2D",X"03",X"2D",X"04",X"2D",X"04",X"2D",X"05",X"2D",X"05",X"2D",X"04",X"12",X"04",X"12",
		X"04",X"11",X"04",X"11",X"05",X"11",X"05",X"11",X"05",X"17",X"05",X"17",X"06",X"17",X"06",X"17",
		X"02",X"3C",X"03",X"3C",X"03",X"3C",X"04",X"3C",X"04",X"3C",X"05",X"3C",X"05",X"19",X"05",X"19",
		X"06",X"19",X"06",X"19",X"02",X"45",X"03",X"45",X"03",X"45",X"04",X"45",X"04",X"45",X"05",X"45",
		X"05",X"2D",X"05",X"2D",X"06",X"2D",X"06",X"2D",X"04",X"27",X"04",X"27",X"05",X"27",X"05",X"27",
		X"06",X"27",X"06",X"27",X"05",X"0D",X"05",X"0D",X"06",X"0D",X"06",X"0D",X"02",X"6D",X"03",X"6C",
		X"03",X"6C",X"04",X"6C",X"04",X"6C",X"05",X"6C",X"06",X"0D",X"06",X"0D",X"06",X"07",X"06",X"07",
		X"06",X"07",X"06",X"07",X"02",X"4E",X"03",X"4E",X"03",X"4E",X"04",X"4E",X"04",X"4E",X"05",X"4E",
		X"06",X"07",X"06",X"07",X"06",X"07",X"06",X"07",X"01",X"54",X"02",X"54",X"06",X"07",X"06",X"07",
		X"06",X"07",X"06",X"07",X"01",X"58",X"02",X"58",X"AF",X"32",X"2D",X"80",X"ED",X"43",X"85",X"81",
		X"C9",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"26",X"7B",X"0A",X"0F",X"0F",X"0F",
		X"5F",X"E6",X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",X"26",X"7D",X"0A",X"77",X"03",X"26",
		X"79",X"CB",X"FD",X"EB",X"60",X"69",X"CF",X"22",X"85",X"81",X"21",X"80",X"93",X"3A",X"42",X"80",
		X"87",X"87",X"87",X"D5",X"EF",X"D1",X"EB",X"72",X"2D",X"73",X"60",X"69",X"01",X"40",X"00",X"ED",
		X"B0",X"3A",X"42",X"80",X"3C",X"FE",X"0C",X"38",X"01",X"AF",X"32",X"42",X"80",X"C9",X"3E",X"31",
		X"32",X"7E",X"7F",X"3C",X"32",X"7C",X"7F",X"AF",X"32",X"2E",X"80",X"ED",X"43",X"85",X"81",X"C9",
		X"3E",X"01",X"32",X"2E",X"80",X"ED",X"43",X"85",X"81",X"C9",X"21",X"1E",X"79",X"36",X"02",X"2C",
		X"36",X"00",X"24",X"36",X"F8",X"24",X"36",X"0E",X"2D",X"36",X"80",X"24",X"36",X"00",X"ED",X"43",
		X"85",X"81",X"AF",X"32",X"2F",X"80",X"21",X"76",X"06",X"11",X"02",X"7F",X"06",X"0F",X"7E",X"12",
		X"1C",X"1C",X"23",X"10",X"F9",X"C9",X"41",X"42",X"43",X"44",X"45",X"46",X"47",X"48",X"49",X"52",
		X"51",X"50",X"4F",X"4A",X"4B",X"ED",X"43",X"85",X"81",X"3E",X"01",X"32",X"2F",X"80",X"C9",X"2A",
		X"85",X"81",X"3A",X"11",X"80",X"BE",X"C0",X"23",X"4D",X"44",X"03",X"7E",X"21",X"A9",X"06",X"D7",
		X"7E",X"21",X"01",X"07",X"CF",X"5E",X"23",X"56",X"EB",X"E9",X"00",X"02",X"03",X"04",X"05",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"0E",X"0E",X"01",X"00",X"01",X"01",X"01",X"01",X"01",X"06",X"07",X"08",X"09",X"01",
		X"01",X"0A",X"0B",X"0C",X"0D",X"01",X"01",X"0F",X"10",X"11",X"00",X"00",X"12",X"13",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"14",X"15",X"16",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"17",X"31",X"07",X"3F",X"07",X"BD",X"03",X"D1",X"03",X"EF",X"03",X"FD",X"03",X"5D",X"07",X"D8",
		X"05",X"3E",X"04",X"48",X"04",X"8E",X"04",X"52",X"04",X"5C",X"04",X"66",X"04",X"67",X"07",X"E1",
		X"05",X"70",X"04",X"7A",X"04",X"2E",X"06",X"40",X"06",X"4A",X"06",X"85",X"06",X"84",X"04",X"0C",
		X"04",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"ED",X"43",X"85",X"81",X"C9",X"26",
		X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",X"26",X"7B",X"0A",X"0F",X"0F",X"0F",X"5F",X"E6",
		X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",X"ED",X"43",X"85",X"81",X"C9",X"0A",X"32",X"22",
		X"84",X"03",X"ED",X"43",X"85",X"81",X"C9",X"26",X"7F",X"0A",X"6F",X"0B",X"0A",X"77",X"03",X"03",
		X"26",X"7B",X"0A",X"0F",X"0F",X"0F",X"5F",X"E6",X"E0",X"77",X"2C",X"7B",X"E6",X"1F",X"77",X"03",
		X"2D",X"26",X"7E",X"0A",X"77",X"03",X"ED",X"43",X"85",X"81",X"C9",X"F7",X"3A",X"11",X"80",X"FE",
		X"0E",X"C8",X"F7",X"3A",X"11",X"80",X"FE",X"0E",X"C0",X"3A",X"87",X"81",X"3C",X"FE",X"10",X"20",
		X"02",X"3E",X"06",X"32",X"87",X"81",X"4F",X"21",X"BD",X"07",X"D7",X"7E",X"32",X"13",X"80",X"79",
		X"21",X"00",X"10",X"CF",X"5E",X"23",X"56",X"ED",X"53",X"85",X"81",X"18",X"CE",X"24",X"00",X"54",
		X"0E",X"40",X"1A",X"64",X"04",X"2A",X"5C",X"0E",X"04",X"38",X"54",X"1A",X"00",X"3A",X"AD",X"85",
		X"FE",X"00",X"C8",X"3A",X"01",X"80",X"0F",X"0F",X"0F",X"0F",X"E6",X"01",X"47",X"21",X"00",X"18",
		X"11",X"00",X"05",X"3A",X"21",X"80",X"A7",X"28",X"01",X"EB",X"4F",X"CD",X"0F",X"08",X"EB",X"3A",
		X"22",X"80",X"A7",X"3E",X"06",X"28",X"07",X"79",X"EE",X"01",X"4F",X"79",X"87",X"81",X"11",X"1F",
		X"08",X"EB",X"D7",X"EB",X"01",X"C0",X"03",X"1A",X"CD",X"28",X"08",X"13",X"10",X"F9",X"C9",X"D5",
		X"C5",X"3A",X"23",X"80",X"A0",X"28",X"02",X"0E",X"02",X"CD",X"FB",X"07",X"C1",X"D1",X"C9",X"01",
		X"1E",X"19",X"02",X"1E",X"19",X"24",X"24",X"24",X"E5",X"F5",X"CD",X"32",X"08",X"F1",X"77",X"E1",
		X"25",X"C9",X"3A",X"03",X"80",X"25",X"A7",X"3E",X"04",X"28",X"03",X"25",X"3E",X"18",X"85",X"E6",
		X"3F",X"6F",X"3E",X"03",X"84",X"0F",X"0F",X"67",X"E6",X"C0",X"B5",X"6F",X"7C",X"E6",X"07",X"81",
		X"67",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"96",
		X"20",X"10",X"C8",X"10",X"AF",X"11",X"3D",X"12",X"CD",X"12",X"A8",X"13",X"73",X"14",X"3F",X"15",
		X"9C",X"16",X"E8",X"16",X"42",X"18",X"24",X"19",X"7A",X"1A",X"29",X"1B",X"77",X"1B",X"F0",X"1C",
		X"0C",X"53",X"00",X"0C",X"FF",X"24",X"0F",X"FF",X"25",X"FF",X"FF",X"28",X"12",X"FF",X"29",X"1F",
		X"FE",X"2A",X"07",X"FE",X"2F",X"1F",X"FE",X"30",X"1F",X"FE",X"2B",X"07",X"FD",X"03",X"EB",X"03",
		X"D7",X"03",X"D6",X"1E",X"04",X"80",X"D6",X"1F",X"06",X"70",X"C3",X"05",X"B7",X"03",X"B6",X"1E",
		X"08",X"80",X"B6",X"26",X"0A",X"70",X"AB",X"1E",X"0C",X"58",X"A9",X"26",X"0E",X"58",X"A1",X"1F",
		X"10",X"40",X"9F",X"26",X"12",X"50",X"9F",X"05",X"9B",X"57",X"9B",X"57",X"93",X"03",X"83",X"03",
		X"7A",X"26",X"14",X"70",X"78",X"1F",X"16",X"70",X"73",X"03",X"69",X"1D",X"18",X"20",X"61",X"2C",
		X"1A",X"5A",X"60",X"25",X"1F",X"5F",X"57",X"5F",X"57",X"5E",X"2C",X"1C",X"5A",X"5B",X"2C",X"1E",
		X"5A",X"5B",X"03",X"53",X"03",X"47",X"03",X"44",X"54",X"00",X"3C",X"1E",X"04",X"60",X"3C",X"26",
		X"06",X"70",X"3B",X"02",X"03",X"27",X"1F",X"08",X"28",X"25",X"26",X"0A",X"38",X"23",X"1F",X"0C",
		X"48",X"23",X"26",X"0E",X"C0",X"21",X"26",X"10",X"58",X"1F",X"1F",X"12",X"68",X"17",X"05",X"17",
		X"1D",X"14",X"D0",X"15",X"2D",X"16",X"68",X"0D",X"FF",X"02",X"01",X"EF",X"05",X"E7",X"2E",X"04",
		X"9C",X"03",X"40",X"00",X"38",X"1C",X"FF",X"18",X"DD",X"26",X"06",X"70",X"DD",X"1E",X"08",X"60",
		X"D3",X"1F",X"0A",X"D0",X"D3",X"26",X"0C",X"C0",X"C9",X"26",X"0E",X"70",X"C9",X"26",X"10",X"60",
		X"C3",X"03",X"BB",X"2E",X"12",X"94",X"03",X"68",X"00",X"20",X"02",X"FF",X"00",X"B3",X"26",X"14",
		X"68",X"B3",X"05",X"A7",X"2E",X"16",X"94",X"03",X"58",X"00",X"C0",X"18",X"FF",X"00",X"A3",X"26",
		X"18",X"70",X"A3",X"1F",X"1A",X"60",X"A3",X"03",X"95",X"26",X"1C",X"68",X"93",X"03",X"83",X"05",
		X"79",X"1F",X"1E",X"D0",X"6F",X"26",X"04",X"70",X"6F",X"1F",X"06",X"60",X"6D",X"1F",X"08",X"70",
		X"6D",X"26",X"0A",X"60",X"67",X"1D",X"0C",X"20",X"67",X"2E",X"0E",X"D8",X"04",X"48",X"1C",X"50",
		X"00",X"20",X"1C",X"FF",X"00",X"5B",X"03",X"4B",X"05",X"47",X"2E",X"10",X"A4",X"04",X"08",X"00",
		X"50",X"08",X"60",X"00",X"C0",X"02",X"44",X"2E",X"12",X"34",X"03",X"78",X"00",X"A8",X"04",X"C0",
		X"06",X"3E",X"1D",X"14",X"70",X"39",X"1F",X"16",X"D0",X"39",X"26",X"18",X"C0",X"33",X"03",X"27",
		X"1E",X"1A",X"90",X"25",X"1F",X"1C",X"80",X"25",X"2E",X"1E",X"60",X"02",X"90",X"04",X"C0",X"08",
		X"23",X"1E",X"04",X"70",X"23",X"05",X"21",X"1F",X"06",X"60",X"1F",X"1E",X"08",X"50",X"1C",X"28",
		X"18",X"1B",X"02",X"01",X"17",X"26",X"0A",X"A0",X"17",X"26",X"0C",X"90",X"15",X"05",X"13",X"1F",
		X"0E",X"B0",X"13",X"1B",X"10",X"A0",X"13",X"1B",X"12",X"90",X"13",X"1F",X"14",X"80",X"0D",X"FF",
		X"22",X"04",X"FF",X"28",X"14",X"EF",X"1F",X"16",X"40",X"E4",X"22",X"02",X"BD",X"26",X"18",X"A0",
		X"BB",X"1F",X"1A",X"A0",X"B8",X"22",X"02",X"A3",X"20",X"1C",X"C0",X"9F",X"1D",X"04",X"E0",X"93",
		X"0F",X"74",X"91",X"26",X"06",X"80",X"8F",X"1E",X"08",X"80",X"8C",X"54",X"00",X"87",X"1E",X"0A",
		X"90",X"87",X"1F",X"0C",X"80",X"83",X"23",X"83",X"57",X"7B",X"03",X"6B",X"1F",X"0E",X"D0",X"6B",
		X"26",X"10",X"A0",X"63",X"05",X"63",X"26",X"12",X"60",X"5B",X"1F",X"14",X"60",X"57",X"36",X"16",
		X"78",X"57",X"03",X"4B",X"57",X"49",X"1F",X"18",X"D0",X"49",X"26",X"1A",X"A0",X"43",X"03",X"36",
		X"1E",X"1C",X"C0",X"36",X"26",X"1E",X"A8",X"36",X"1F",X"04",X"90",X"36",X"1E",X"06",X"78",X"2C",
		X"1F",X"08",X"90",X"2B",X"05",X"1F",X"1F",X"0A",X"80",X"1F",X"26",X"0C",X"60",X"1F",X"1F",X"0E",
		X"40",X"18",X"24",X"03",X"17",X"21",X"10",X"60",X"17",X"1D",X"14",X"20",X"0D",X"FF",X"02",X"01",
		X"F0",X"05",X"ED",X"2E",X"16",X"9C",X"03",X"A0",X"00",X"80",X"10",X"80",X"00",X"E3",X"2E",X"18",
		X"2C",X"02",X"90",X"00",X"80",X"1C",X"DB",X"1E",X"1A",X"60",X"DB",X"1F",X"1C",X"50",X"D1",X"2E",
		X"1E",X"7C",X"03",X"38",X"00",X"80",X"02",X"C0",X"00",X"CB",X"03",X"C5",X"26",X"04",X"B0",X"C5",
		X"1F",X"06",X"A0",X"C5",X"1D",X"08",X"60",X"BD",X"2E",X"0A",X"24",X"03",X"48",X"00",X"28",X"02",
		X"FF",X"00",X"BB",X"05",X"AF",X"1F",X"0C",X"50",X"AD",X"1F",X"0E",X"40",X"AA",X"26",X"10",X"50",
		X"A7",X"26",X"12",X"40",X"A7",X"2E",X"14",X"24",X"04",X"60",X"00",X"D8",X"10",X"28",X"08",X"FF",
		X"02",X"9F",X"03",X"8B",X"05",X"87",X"22",X"01",X"83",X"23",X"73",X"02",X"45",X"73",X"4E",X"2F",
		X"73",X"4C",X"63",X"05",X"5F",X"02",X"45",X"4F",X"05",X"3F",X"22",X"04",X"33",X"23",X"31",X"23",
		X"2B",X"23",X"2B",X"57",X"28",X"03",X"20",X"4D",X"20",X"03",X"10",X"03",X"0D",X"FF",X"24",X"07",
		X"FF",X"2F",X"0F",X"FE",X"30",X"0F",X"FE",X"28",X"1C",X"FD",X"03",X"EF",X"03",X"E3",X"57",X"E3",
		X"05",X"DD",X"1F",X"04",X"A0",X"DD",X"1E",X"06",X"90",X"DB",X"21",X"08",X"70",X"DB",X"1E",X"0C",
		X"A0",X"DB",X"1F",X"0E",X"90",X"D1",X"3D",X"10",X"C0",X"CB",X"03",X"BF",X"3E",X"12",X"A0",X"BB",
		X"03",X"BB",X"3E",X"14",X"60",X"B7",X"3E",X"16",X"A0",X"B3",X"03",X"B3",X"3F",X"18",X"60",X"AF",
		X"3F",X"1A",X"20",X"A7",X"05",X"A5",X"21",X"1C",X"68",X"9B",X"3E",X"04",X"40",X"97",X"3E",X"06",
		X"80",X"95",X"3E",X"08",X"A0",X"93",X"3E",X"0A",X"C0",X"93",X"03",X"7B",X"05",X"7B",X"54",X"00",
		X"71",X"2E",X"0C",X"60",X"0C",X"30",X"00",X"30",X"10",X"30",X"18",X"30",X"08",X"30",X"00",X"30",
		X"10",X"30",X"18",X"30",X"08",X"30",X"00",X"30",X"10",X"30",X"18",X"30",X"08",X"71",X"1D",X"0E",
		X"20",X"70",X"25",X"0F",X"70",X"24",X"0F",X"6B",X"1E",X"10",X"80",X"69",X"26",X"12",X"80",X"67",
		X"1E",X"14",X"80",X"65",X"26",X"16",X"80",X"63",X"03",X"4B",X"05",X"4B",X"1F",X"18",X"C0",X"3F",
		X"03",X"35",X"1F",X"1A",X"80",X"32",X"2E",X"1C",X"D8",X"03",X"C0",X"18",X"18",X"10",X"C0",X"08",
		X"31",X"1D",X"1E",X"40",X"2F",X"05",X"23",X"2E",X"04",X"C0",X"01",X"C0",X"18",X"20",X"2E",X"06",
		X"20",X"01",X"C0",X"08",X"1D",X"2E",X"08",X"C0",X"01",X"C0",X"18",X"17",X"1F",X"0A",X"C0",X"17",
		X"21",X"0C",X"80",X"17",X"1F",X"10",X"40",X"0D",X"FF",X"24",X"07",X"F3",X"26",X"04",X"C0",X"F3",
		X"1E",X"06",X"B0",X"EB",X"2E",X"08",X"3C",X"03",X"C0",X"00",X"C0",X"10",X"C0",X"00",X"DB",X"2E",
		X"0A",X"34",X"02",X"20",X"02",X"FF",X"00",X"D7",X"1F",X"0C",X"C0",X"D5",X"26",X"0E",X"D0",X"D5",
		X"30",X"FF",X"CB",X"2E",X"10",X"1C",X"03",X"98",X"00",X"80",X"02",X"40",X"00",X"BB",X"2E",X"12",
		X"1C",X"01",X"FF",X"00",X"B6",X"1E",X"14",X"C0",X"B6",X"26",X"16",X"D0",X"B4",X"30",X"0F",X"AA",
		X"1F",X"18",X"B0",X"AA",X"1F",X"1A",X"A0",X"9F",X"21",X"1C",X"A0",X"9B",X"03",X"8B",X"1D",X"04",
		X"30",X"83",X"05",X"77",X"2D",X"06",X"C0",X"6F",X"3A",X"10",X"48",X"6B",X"38",X"12",X"60",X"6B",
		X"38",X"14",X"30",X"67",X"38",X"16",X"48",X"5F",X"1F",X"18",X"80",X"5D",X"26",X"1A",X"70",X"56",
		X"2E",X"1C",X"14",X"0B",X"40",X"00",X"38",X"04",X"50",X"06",X"38",X"04",X"3C",X"08",X"30",X"04",
		X"20",X"00",X"20",X"10",X"20",X"00",X"20",X"10",X"20",X"00",X"55",X"26",X"1E",X"70",X"4F",X"26",
		X"04",X"80",X"4F",X"1D",X"06",X"D0",X"48",X"2E",X"08",X"D8",X"03",X"08",X"00",X"58",X"18",X"FF",
		X"00",X"41",X"2E",X"0A",X"48",X"02",X"78",X"00",X"FF",X"08",X"33",X"1F",X"0C",X"70",X"27",X"26",
		X"0E",X"70",X"25",X"26",X"10",X"90",X"23",X"26",X"12",X"B0",X"17",X"21",X"14",X"C0",X"17",X"21",
		X"18",X"A0",X"0D",X"FF",X"22",X"08",X"F1",X"1F",X"04",X"80",X"EF",X"1E",X"06",X"80",X"ED",X"22",
		X"03",X"CA",X"30",X"3F",X"C9",X"2E",X"08",X"70",X"06",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",
		X"1C",X"60",X"00",X"60",X"04",X"C6",X"2E",X"0A",X"58",X"06",X"30",X"04",X"60",X"0C",X"60",X"10",
		X"60",X"14",X"60",X"1C",X"60",X"00",X"C3",X"2E",X"0C",X"40",X"06",X"60",X"04",X"60",X"0C",X"60",
		X"10",X"60",X"14",X"60",X"1C",X"60",X"00",X"C0",X"2E",X"0E",X"40",X"06",X"30",X"00",X"60",X"04",
		X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"BD",X"2E",X"10",X"40",X"06",X"60",X"00",X"60",
		X"04",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"BA",X"2E",X"12",X"58",X"07",X"30",X"1C",
		X"60",X"00",X"60",X"04",X"60",X"0C",X"60",X"10",X"60",X"14",X"60",X"1C",X"A7",X"2F",X"07",X"A1",
		X"1E",X"14",X"70",X"9F",X"26",X"16",X"60",X"9E",X"22",X"02",X"9D",X"1F",X"18",X"50",X"9B",X"1E",
		X"1A",X"40",X"83",X"10",X"74",X"81",X"26",X"1C",X"40",X"7B",X"1D",X"1E",X"D8",X"6C",X"23",X"6B",
		X"1E",X"04",X"B0",X"6B",X"1F",X"06",X"80",X"6B",X"1E",X"08",X"50",X"6B",X"1F",X"0A",X"20",X"66",
		X"54",X"00",X"4F",X"22",X"10",X"36",X"1F",X"0C",X"48",X"36",X"1F",X"0E",X"20",X"2B",X"3B",X"10",
		X"C0",X"27",X"3C",X"12",X"A0",X"17",X"11",X"76",X"11",X"1D",X"14",X"20",X"0F",X"23",X"0D",X"F3",
		X"03",X"F3",X"30",X"FF",X"F3",X"57",X"EE",X"2E",X"04",X"14",X"05",X"08",X"00",X"A0",X"08",X"30",
		X"0C",X"FF",X"10",X"FF",X"00",X"EA",X"05",X"E5",X"26",X"06",X"30",X"E5",X"26",X"08",X"C8",X"E2",
		X"1F",X"0A",X"48",X"E2",X"1F",X"0C",X"B0",X"DF",X"26",X"0E",X"60",X"DF",X"26",X"10",X"98",X"CC",
		X"1E",X"12",X"40",X"C8",X"26",X"14",X"60",X"C8",X"26",X"16",X"20",X"C7",X"21",X"18",X"48",X"C3",
		X"1E",X"1C",X"40",X"BB",X"57",X"B3",X"1F",X"1E",X"48",X"A8",X"03",X"A5",X"2E",X"04",X"A0",X"02",
		X"B0",X"02",X"80",X"00",X"A5",X"2E",X"06",X"74",X"04",X"78",X"00",X"50",X"18",X"50",X"08",X"80",
		X"00",X"A5",X"2E",X"08",X"14",X"04",X"78",X"00",X"50",X"08",X"50",X"18",X"80",X"00",X"9B",X"05",
		X"93",X"2E",X"0A",X"7C",X"05",X"A0",X"00",X"F0",X"10",X"30",X"0F",X"30",X"1F",X"80",X"00",X"93",
		X"1F",X"0C",X"50",X"93",X"26",X"0E",X"40",X"93",X"2E",X"10",X"14",X"03",X"AC",X"00",X"FF",X"10",
		X"80",X"00",X"83",X"03",X"7F",X"2E",X"12",X"84",X"07",X"50",X"00",X"C0",X"10",X"50",X"10",X"28",
		X"0B",X"50",X"10",X"70",X"0C",X"60",X"0D",X"77",X"1D",X"14",X"D0",X"73",X"05",X"73",X"26",X"04",
		X"58",X"73",X"1F",X"06",X"48",X"6D",X"2E",X"16",X"14",X"01",X"80",X"00",X"6A",X"2E",X"18",X"14",
		X"01",X"80",X"00",X"67",X"2E",X"1A",X"14",X"01",X"80",X"00",X"64",X"35",X"1C",X"14",X"61",X"35",
		X"1E",X"14",X"47",X"2E",X"08",X"80",X"06",X"08",X"00",X"58",X"08",X"60",X"00",X"60",X"02",X"80",
		X"00",X"60",X"04",X"47",X"2E",X"0A",X"68",X"08",X"08",X"00",X"88",X"08",X"60",X"00",X"60",X"1C",
		X"38",X"00",X"18",X"12",X"A8",X"14",X"80",X"00",X"47",X"2E",X"0C",X"50",X"03",X"08",X"00",X"78",
		X"18",X"80",X"00",X"37",X"1B",X"0E",X"B8",X"37",X"1B",X"10",X"48",X"27",X"2E",X"12",X"50",X"02",
		X"68",X"04",X"E0",X"08",X"24",X"2E",X"14",X"38",X"02",X"98",X"04",X"E0",X"08",X"21",X"2E",X"16",
		X"20",X"02",X"C8",X"04",X"E0",X"08",X"1F",X"2E",X"18",X"90",X"03",X"08",X"1C",X"E0",X"00",X"D0",
		X"08",X"1C",X"2E",X"1A",X"A8",X"03",X"38",X"1C",X"E0",X"00",X"D0",X"08",X"19",X"2E",X"1C",X"C0",
		X"03",X"68",X"1C",X"E0",X"00",X"D0",X"08",X"19",X"1F",X"1E",X"88",X"19",X"1F",X"04",X"68",X"19",
		X"1F",X"06",X"48",X"13",X"1B",X"08",X"88",X"13",X"1B",X"0C",X"48",X"0D",X"FB",X"02",X"1F",X"F5",
		X"1D",X"10",X"A0",X"F3",X"1D",X"12",X"80",X"F1",X"1D",X"14",X"60",X"EF",X"1D",X"16",X"40",X"EB",
		X"05",X"E3",X"02",X"38",X"D5",X"21",X"18",X"50",X"D3",X"05",X"D1",X"57",X"CF",X"03",X"C7",X"03",
		X"C3",X"02",X"6F",X"BF",X"05",X"B3",X"33",X"9F",X"34",X"87",X"18",X"76",X"85",X"4E",X"0F",X"83",
		X"4C",X"73",X"02",X"45",X"63",X"05",X"63",X"57",X"5B",X"02",X"65",X"4B",X"05",X"3F",X"03",X"2F",
		X"03",X"20",X"4D",X"1F",X"03",X"10",X"05",X"0D",X"FF",X"03",X"FF",X"30",X"3F",X"F7",X"05",X"F3",
		X"57",X"EF",X"03",X"E3",X"05",X"DB",X"03",X"CF",X"05",X"C6",X"2E",X"1C",X"D8",X"08",X"60",X"14",
		X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"C6",X"2E",
		X"1E",X"98",X"08",X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"60",
		X"10",X"60",X"00",X"C6",X"2E",X"04",X"58",X"08",X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",X"1C",
		X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",X"1C",X"BE",X"2E",X"06",X"B8",X"08",X"40",X"08",X"60",
		X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"BE",X"2E",X"08",
		X"78",X"08",X"40",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",X"60",X"08",X"60",X"18",
		X"60",X"08",X"B8",X"2E",X"0A",X"C8",X"07",X"40",X"1C",X"60",X"0C",X"60",X"1C",X"60",X"0C",X"60",
		X"1C",X"60",X"0C",X"60",X"1C",X"B8",X"2E",X"0C",X"98",X"07",X"40",X"00",X"60",X"10",X"60",X"00",
		X"60",X"10",X"60",X"00",X"60",X"10",X"60",X"00",X"B8",X"2E",X"0E",X"68",X"07",X"40",X"04",X"60",
		X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"60",X"14",X"60",X"04",X"A9",X"1E",X"10",X"B0",X"A9",
		X"1E",X"12",X"90",X"A7",X"1E",X"14",X"A0",X"A5",X"1E",X"16",X"B0",X"A5",X"1E",X"18",X"90",X"9B",
		X"18",X"76",X"91",X"1F",X"1A",X"40",X"8F",X"1F",X"1C",X"40",X"8B",X"18",X"76",X"87",X"1E",X"1E",
		X"50",X"87",X"1E",X"04",X"40",X"7B",X"18",X"76",X"6F",X"1F",X"06",X"C0",X"6F",X"1E",X"08",X"A0",
		X"6F",X"1F",X"0A",X"80",X"64",X"2E",X"0C",X"98",X"10",X"80",X"18",X"80",X"10",X"80",X"09",X"20",
		X"0C",X"40",X"18",X"20",X"1A",X"10",X"18",X"28",X"10",X"10",X"08",X"20",X"06",X"48",X"08",X"18",
		X"0C",X"70",X"18",X"A0",X"13",X"98",X"08",X"80",X"04",X"47",X"1D",X"0E",X"C0",X"47",X"1D",X"10",
		X"A0",X"47",X"1D",X"12",X"80",X"47",X"1D",X"14",X"60",X"43",X"1D",X"16",X"C0",X"43",X"1D",X"18",
		X"A0",X"43",X"1D",X"1A",X"80",X"43",X"1D",X"1C",X"60",X"36",X"1E",X"1E",X"80",X"36",X"26",X"04",
		X"60",X"36",X"1E",X"06",X"40",X"2B",X"1F",X"08",X"50",X"21",X"20",X"0A",X"80",X"1B",X"20",X"0E",
		X"80",X"19",X"1B",X"12",X"D0",X"19",X"1B",X"14",X"20",X"13",X"1B",X"16",X"D0",X"13",X"1B",X"18",
		X"20",X"0D",X"FB",X"11",X"74",X"F3",X"22",X"08",X"E9",X"2D",X"04",X"60",X"E6",X"22",X"08",X"E4",
		X"2E",X"0E",X"9C",X"01",X"80",X"00",X"DC",X"2E",X"10",X"2C",X"02",X"F8",X"00",X"40",X"1C",X"CB",
		X"26",X"12",X"B0",X"CB",X"1F",X"14",X"A0",X"CB",X"2E",X"16",X"2C",X"07",X"70",X"00",X"E8",X"10",
		X"20",X"12",X"B8",X"10",X"B8",X"00",X"20",X"02",X"20",X"00",X"C3",X"23",X"C3",X"35",X"18",X"7C",
		X"BF",X"35",X"1A",X"7C",X"BB",X"35",X"1C",X"7C",X"B7",X"39",X"1E",X"7C",X"AF",X"3B",X"04",X"24",
		X"A7",X"3B",X"06",X"24",X"A3",X"22",X"0C",X"9B",X"03",X"8B",X"05",X"8B",X"1D",X"08",X"70",X"84",
		X"1D",X"0A",X"70",X"84",X"22",X"04",X"77",X"2E",X"0C",X"34",X"09",X"60",X"00",X"A0",X"10",X"28",
		X"0D",X"50",X"10",X"70",X"0C",X"60",X"0D",X"40",X"06",X"30",X"04",X"20",X"08",X"75",X"1F",X"0E",
		X"60",X"73",X"1E",X"10",X"70",X"73",X"23",X"71",X"1F",X"12",X"80",X"6F",X"1E",X"14",X"90",X"6D",
		X"1F",X"16",X"A0",X"6B",X"1E",X"18",X"B0",X"69",X"1F",X"1A",X"C0",X"67",X"1E",X"1C",X"D0",X"67",
		X"57",X"63",X"03",X"63",X"03",X"53",X"22",X"10",X"43",X"03",X"3B",X"05",X"2B",X"2E",X"1E",X"E0",
		X"05",X"08",X"00",X"60",X"18",X"20",X"1C",X"D8",X"18",X"20",X"14",X"27",X"21",X"04",X"68",X"23",
		X"23",X"1E",X"1D",X"08",X"20",X"1D",X"1F",X"0A",X"D0",X"1D",X"1F",X"0C",X"A0",X"1B",X"1D",X"0E",
		X"38",X"18",X"1D",X"10",X"50",X"17",X"1E",X"12",X"D0",X"17",X"1E",X"14",X"A0",X"15",X"1D",X"16",
		X"68",X"13",X"23",X"0D",X"FF",X"30",X"0F",X"FF",X"29",X"0F",X"FF",X"2B",X"03",X"FF",X"2A",X"03",
		X"F3",X"57",X"EE",X"2E",X"04",X"14",X"09",X"08",X"00",X"A0",X"08",X"30",X"0C",X"48",X"10",X"30",
		X"00",X"50",X"10",X"68",X"00",X"30",X"1C",X"20",X"18",X"E5",X"1B",X"06",X"C0",X"E5",X"1F",X"08",
		X"B0",X"E5",X"1F",X"0A",X"48",X"E5",X"1B",X"0C",X"38",X"E3",X"1F",X"0E",X"C0",X"E3",X"1B",X"10",
		X"B0",X"E3",X"1B",X"12",X"48",X"E3",X"1F",X"14",X"38",X"DC",X"2E",X"16",X"7C",X"04",X"08",X"10",
		X"78",X"00",X"50",X"10",X"40",X"00",X"C9",X"35",X"18",X"48",X"C9",X"35",X"1A",X"38",X"C7",X"35",
		X"1C",X"48",X"C7",X"35",X"1E",X"38",X"BD",X"1E",X"04",X"B0",X"BB",X"1E",X"06",X"B0",X"BB",X"1E",
		X"08",X"90",X"B9",X"1E",X"0A",X"90",X"B3",X"2E",X"0C",X"CC",X"01",X"20",X"00",X"A7",X"2E",X"0E",
		X"74",X"04",X"58",X"00",X"A0",X"18",X"A0",X"08",X"20",X"00",X"A3",X"2E",X"10",X"14",X"01",X"20",
		X"00",X"A3",X"57",X"A1",X"2E",X"12",X"14",X"01",X"20",X"00",X"97",X"03",X"93",X"2E",X"14",X"7C",
		X"02",X"98",X"00",X"20",X"02",X"8D",X"1D",X"16",X"E0",X"8D",X"1D",X"18",X"D0",X"8B",X"1D",X"1A",
		X"E0",X"8B",X"1D",X"1C",X"D0",X"87",X"05",X"83",X"03",X"77",X"1E",X"1E",X"60",X"77",X"1F",X"04",
		X"50",X"73",X"05",X"73",X"2E",X"06",X"14",X"04",X"70",X"00",X"E0",X"10",X"A0",X"10",X"20",X"00",
		X"6F",X"1F",X"08",X"60",X"6F",X"1E",X"0A",X"50",X"6B",X"03",X"5B",X"05",X"55",X"1B",X"0C",X"A8",
		X"47",X"2E",X"0E",X"78",X"03",X"08",X"00",X"C8",X"18",X"20",X"00",X"47",X"2E",X"10",X"90",X"03",
		X"08",X"00",X"F8",X"18",X"20",X"00",X"47",X"2E",X"12",X"A8",X"04",X"08",X"00",X"E0",X"18",X"48",
		X"18",X"20",X"00",X"37",X"1F",X"14",X"C0",X"37",X"1F",X"16",X"B0",X"30",X"1B",X"18",X"68",X"2E",
		X"1B",X"1A",X"58",X"2C",X"1B",X"1C",X"48",X"2A",X"1B",X"1E",X"38",X"27",X"36",X"04",X"14",X"23",
		X"36",X"06",X"14",X"1F",X"36",X"08",X"14",X"1B",X"39",X"0A",X"14",X"18",X"2E",X"0C",X"88",X"08",
		X"40",X"00",X"80",X"18",X"80",X"10",X"80",X"08",X"80",X"00",X"80",X"18",X"80",X"10",X"80",X"08",
		X"18",X"2E",X"0E",X"48",X"08",X"40",X"10",X"80",X"08",X"80",X"00",X"80",X"18",X"80",X"10",X"80",
		X"08",X"80",X"00",X"80",X"18",X"17",X"21",X"10",X"70",X"0D",X"F7",X"1B",X"14",X"20",X"F3",X"1B",
		X"16",X"A0",X"F3",X"1B",X"18",X"70",X"ED",X"1F",X"1A",X"A0",X"EB",X"1F",X"1C",X"90",X"E9",X"1F",
		X"1E",X"80",X"E7",X"1F",X"04",X"70",X"E3",X"57",X"DF",X"1B",X"06",X"C0",X"D9",X"1B",X"08",X"C0",
		X"D3",X"03",X"BB",X"05",X"B1",X"21",X"0A",X"B0",X"B1",X"21",X"0E",X"50",X"AB",X"03",X"A1",X"3E",
		X"12",X"90",X"9D",X"3E",X"14",X"70",X"99",X"40",X"16",X"50",X"95",X"3E",X"18",X"30",X"93",X"05",
		X"8D",X"40",X"1A",X"50",X"89",X"3E",X"1C",X"70",X"85",X"3E",X"1E",X"90",X"81",X"3E",X"04",X"B0",
		X"7B",X"03",X"71",X"1F",X"06",X"D0",X"6F",X"26",X"08",X"C0",X"6D",X"1F",X"0A",X"B0",X"6B",X"26",
		X"0C",X"A0",X"69",X"1F",X"0E",X"90",X"63",X"05",X"5F",X"57",X"5B",X"02",X"EC",X"43",X"05",X"40",
		X"1D",X"10",X"30",X"40",X"1D",X"12",X"20",X"3B",X"03",X"36",X"1B",X"14",X"C0",X"25",X"2E",X"16",
		X"E0",X"02",X"C0",X"18",X"C0",X"08",X"25",X"2E",X"18",X"10",X"02",X"C0",X"08",X"C0",X"18",X"23",
		X"2E",X"1A",X"D0",X"02",X"A0",X"18",X"A0",X"08",X"23",X"2E",X"1C",X"20",X"02",X"A0",X"08",X"A0",
		X"18",X"23",X"05",X"1B",X"02",X"E6",X"0E",X"05",X"0D",X"FF",X"02",X"6D",X"F7",X"05",X"F3",X"22",
		X"02",X"E7",X"23",X"E7",X"4E",X"0F",X"E7",X"02",X"F1",X"E3",X"4C",X"DF",X"05",X"DB",X"02",X"34",
		X"D5",X"05",X"CB",X"02",X"49",X"C5",X"05",X"BB",X"02",X"3E",X"BB",X"4D",X"AB",X"05",X"A1",X"33",
		X"8F",X"34",X"7F",X"02",X"46",X"77",X"05",X"73",X"18",X"76",X"67",X"4C",X"67",X"02",X"66",X"65",
		X"05",X"5B",X"02",X"21",X"55",X"05",X"4B",X"03",X"3B",X"05",X"37",X"57",X"33",X"4D",X"33",X"03",
		X"23",X"05",X"1B",X"03",X"1F",X"05",X"0D",X"FF",X"02",X"08",X"F3",X"05",X"EF",X"2E",X"04",X"3C",
		X"05",X"80",X"00",X"80",X"10",X"70",X"00",X"70",X"10",X"70",X"00",X"EE",X"1D",X"06",X"D0",X"EE",
		X"26",X"08",X"80",X"E6",X"2E",X"0A",X"3C",X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"E5",X"1F",
		X"0C",X"80",X"DE",X"2E",X"0E",X"3C",X"03",X"60",X"00",X"60",X"10",X"60",X"00",X"D7",X"1F",X"10",
		X"C0",X"D7",X"2E",X"12",X"26",X"06",X"50",X"02",X"78",X"12",X"18",X"10",X"18",X"00",X"80",X"02",
		X"20",X"00",X"D5",X"1F",X"14",X"D0",X"D2",X"26",X"16",X"50",X"CD",X"2E",X"18",X"1C",X"04",X"40",
		X"00",X"A0",X"10",X"D8",X"00",X"20",X"02",X"C6",X"1F",X"04",X"50",X"C2",X"2E",X"1A",X"1C",X"03",
		X"80",X"00",X"A0",X"00",X"20",X"02",X"BE",X"35",X"1C",X"1C",X"BA",X"3B",X"1E",X"1C",X"B6",X"1F",
		X"06",X"D0",X"B6",X"26",X"08",X"C0",X"B6",X"1D",X"0A",X"50",X"B3",X"03",X"A9",X"1D",X"0C",X"B0",
		X"A3",X"03",X"A0",X"26",X"0E",X"A0",X"A0",X"1F",X"10",X"90",X"93",X"05",X"8B",X"03",X"7B",X"05",
		X"78",X"21",X"12",X"C8",X"76",X"2E",X"16",X"78",X"08",X"50",X"14",X"50",X"04",X"50",X"14",X"50",
		X"04",X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"76",X"2E",X"18",X"18",X"08",X"50",X"0C",
		X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"6B",X"2E",
		X"1A",X"70",X"09",X"40",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",X"1C",X"50",X"0C",X"50",
		X"1C",X"50",X"0C",X"50",X"1C",X"6B",X"2E",X"1C",X"20",X"09",X"40",X"04",X"50",X"14",X"50",X"04",
		X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"50",X"14",X"50",X"04",X"61",X"2E",X"1E",X"A4",
		X"07",X"18",X"00",X"10",X"1C",X"60",X"18",X"38",X"14",X"40",X"16",X"60",X"1E",X"20",X"1C",X"5F",
		X"1F",X"04",X"80",X"5B",X"26",X"06",X"60",X"5B",X"1D",X"08",X"20",X"57",X"1F",X"0A",X"40",X"4E",
		X"2E",X"14",X"AC",X"06",X"50",X"00",X"A8",X"10",X"10",X"08",X"E0",X"18",X"A0",X"10",X"C0",X"00",
		X"48",X"2E",X"12",X"D4",X"06",X"08",X"00",X"90",X"18",X"10",X"08",X"A0",X"18",X"E0",X"10",X"C0",
		X"00",X"47",X"2E",X"10",X"44",X"06",X"18",X"00",X"70",X"08",X"70",X"18",X"C0",X"10",X"F0",X"10",
		X"20",X"18",X"3B",X"26",X"16",X"B0",X"37",X"1F",X"18",X"90",X"1F",X"1B",X"1A",X"90",X"1F",X"1B",
		X"1C",X"70",X"1F",X"1B",X"1E",X"50",X"1B",X"1B",X"04",X"70",X"1B",X"35",X"06",X"24",X"1B",X"02",
		X"3F",X"17",X"3B",X"08",X"24",X"15",X"21",X"0A",X"C0",X"13",X"3B",X"0E",X"24",X"0F",X"05",X"0D",
		X"01",X"57",X"FF",X"03",X"F3",X"1D",X"14",X"20",X"EF",X"05",X"E7",X"2E",X"16",X"9C",X"03",X"40",
		X"00",X"38",X"1C",X"40",X"18",X"E5",X"1B",X"18",X"60",X"E1",X"2E",X"1A",X"24",X"03",X"80",X"00",
		X"80",X"10",X"80",X"00",X"DD",X"2E",X"1C",X"9C",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"D7",
		X"1B",X"1E",X"78",X"D7",X"1B",X"04",X"48",X"D7",X"2E",X"06",X"24",X"03",X"80",X"00",X"80",X"10",
		X"80",X"00",X"D3",X"2E",X"08",X"9C",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"D3",X"1B",X"0A",
		X"60",X"CD",X"2E",X"0C",X"24",X"03",X"80",X"00",X"80",X"10",X"80",X"00",X"CB",X"26",X"0E",X"C8",
		X"CB",X"26",X"10",X"60",X"C5",X"2E",X"12",X"9C",X"08",X"60",X"00",X"78",X"10",X"20",X"12",X"F8",
		X"10",X"58",X"10",X"50",X"18",X"50",X"08",X"20",X"00",X"C5",X"2E",X"14",X"24",X"08",X"60",X"00",
		X"90",X"10",X"20",X"0C",X"E0",X"10",X"58",X"10",X"50",X"08",X"50",X"18",X"20",X"00",X"C5",X"57",
		X"C3",X"03",X"BB",X"3B",X"16",X"70",X"BB",X"3B",X"18",X"50",X"B7",X"3C",X"1A",X"70",X"B7",X"3B",
		X"1C",X"50",X"B3",X"03",X"A3",X"03",X"95",X"1F",X"1E",X"80",X"93",X"05",X"93",X"1F",X"04",X"70",
		X"91",X"1F",X"06",X"60",X"8F",X"1F",X"08",X"50",X"85",X"03",X"7D",X"26",X"0A",X"E0",X"7D",X"26",
		X"0C",X"88",X"7D",X"26",X"0E",X"50",X"79",X"26",X"10",X"C0",X"79",X"26",X"12",X"6C",X"79",X"26",
		X"14",X"18",X"6F",X"21",X"16",X"80",X"6F",X"3B",X"1A",X"34",X"6B",X"3B",X"1C",X"34",X"6B",X"05",
		X"67",X"1D",X"1E",X"B0",X"65",X"1D",X"04",X"A0",X"63",X"03",X"53",X"05",X"4F",X"26",X"06",X"80",
		X"4C",X"1F",X"08",X"68",X"4B",X"2E",X"0A",X"34",X"02",X"A0",X"04",X"20",X"06",X"44",X"1B",X"0C",
		X"70",X"3E",X"1B",X"0E",X"C0",X"3E",X"1D",X"10",X"70",X"3E",X"1B",X"12",X"18",X"38",X"1B",X"14",
		X"70",X"37",X"2E",X"16",X"A4",X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"37",X"2E",X"04",X"34",
		X"03",X"70",X"00",X"70",X"10",X"70",X"00",X"33",X"02",X"E6",X"23",X"05",X"22",X"2E",X"06",X"48",
		X"02",X"B8",X"04",X"20",X"08",X"22",X"2E",X"08",X"34",X"01",X"20",X"00",X"1B",X"2E",X"0A",X"48",
		X"08",X"30",X"00",X"A0",X"04",X"A0",X"10",X"80",X"0C",X"40",X"10",X"80",X"18",X"A0",X"18",X"20",
		X"00",X"17",X"21",X"18",X"90",X"17",X"21",X"1C",X"70",X"17",X"02",X"7E",X"0F",X"05",X"0F",X"30",
		X"1F",X"0D",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"68");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
